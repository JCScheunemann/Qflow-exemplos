* SPICE3 file created from multiplicador.ext - technology: scmos

.option scale=0.05u

C0 B<1> gnd 3.54fF
C1 A<3> gnd 2.85fF
C2 INVX4_4/Y INVX4_1/Y 2.08fF
C3 BUFX4_2/Y vdd 3.57fF
C4 INVX4_3/Y gnd 2.45fF
C5 vdd clk 4.83fF
C6 B<0> vdd 2.70fF
C7 A<4> B<0> 2.05fF
C8 NAND2X1_33/Y gnd 3.31fF
C9 vdd NAND3X1_79/Y 2.08fF
C10 B<5> vdd 3.03fF
C11 NOR3X1_1/C gnd 19.66fF
C12 INVX4_4/Y vdd 3.06fF
C13 AOI21X1_4/B vdd 3.81fF
C14 AOI21X1_7/B INVX1_48/Y 2.18fF
C15 AOI22X1_10/D gnd 4.92fF
C16 INVX1_16/A gnd 3.35fF
C17 XOR2X1_3/Y gnd 4.12fF
C18 B<4> gnd 37.80fF
C19 OAI21X1_7/Y gnd 3.25fF
C20 XOR2X1_1/A gnd 12.56fF
C21 NOR2X1_9/A gnd 5.31fF
C22 INVX2_9/Y vdd 5.46fF
C23 NAND2X1_15/Y gnd 8.26fF
C24 INVX4_6/Y vdd 2.23fF
C25 AND2X2_14/Y gnd 15.12fF
C26 AOI22X1_6/C BUFX2_11/A 2.26fF
C27 AND2X2_18/Y vdd 2.69fF
C28 NAND3X1_25/Y NAND3X1_49/C 2.09fF
C29 NOR3X1_2/C vdd 2.15fF
C30 AND2X2_5/A vdd 2.62fF
C31 NAND3X1_18/B vdd 2.13fF
C32 NOR2X1_35/B vdd 2.24fF
C33 BUFX4_3/Y vdd 4.05fF
C34 AOI21X1_81/B vdd 2.25fF
C35 INVX1_13/A BUFX2_11/A 2.23fF
C36 NAND3X1_91/Y vdd 2.18fF
C37 NAND3X1_22/C vdd 2.37fF
C38 A<2> vdd 4.40fF
C39 INVX2_8/A vdd 2.34fF
C40 INVX4_1/Y vdd 6.34fF
C41 AOI21X1_75/B vdd 2.43fF
C42 B<3> gnd 2.21fF
C43 XOR2X1_4/B gnd 30.22fF
C44 BUFX4_4/A vdd 2.34fF
C45 AOI22X1_6/C AOI22X1_6/D 2.22fF
C46 INVX1_13/Y gnd 69.26fF
C47 INVX1_18/A vdd 2.89fF
C48 INVX2_3/Y vdd 2.54fF
C49 A<5> vdd 2.95fF
C50 vdd NAND3X1_27/C 2.03fF
C51 INVX4_3/Y INVX2_9/Y 3.24fF
C52 XNOR2X1_8/Y XNOR2X1_8/B 2.18fF
C53 OR2X2_1/A vdd 2.33fF
C54 A<6> vdd 2.44fF
C55 BUFX4_2/Y gnd 2.81fF
C56 A<4> vdd 2.20fF
C57 gnd clk 18.89fF
C58 B<0> gnd 3.05fF
C59 AOI21X1_40/Y XNOR2X1_1/Y 2.69fF
C60 INVX1_9/A AOI22X1_6/C 2.34fF
C61 B<5> gnd 19.99fF
C62 NOR2X1_6/Y gnd 2.13fF
C63 AOI22X1_20/A vdd 2.39fF
C64 NAND2X1_85/Y vdd 2.38fF
C65 NOR2X1_4/A gnd 27.89fF
C66 INVX2_1/Y vdd 2.79fF
C67 INVX1_6/Y NAND3X1_27/C 2.01fF
C68 B<1> A<5> 2.18fF
C69 A<1> vdd 2.70fF
C70 OAI21X1_83/Y vdd 2.22fF
C71 A<6> B<1> 2.28fF
C72 AND2X2_18/Y gnd 19.40fF
C73 vdd AOI21X1_78/C 2.16fF
C74 INVX1_9/A BUFX2_11/A 3.20fF
C75 AND2X2_12/Y vdd 2.26fF
C76 BUFX4_1/Y vdd 2.51fF
C77 BUFX4_3/Y gnd 2.12fF
C78 A<3> vdd 4.57fF
C79 B<4> A<2> 3.11fF
C80 gnd INVX1_6/A 2.31fF
C81 AOI21X1_81/C vdd 2.28fF
C82 INVX4_3/Y vdd 6.03fF
C83 NAND3X1_22/C gnd 2.15fF
C84 OAI21X1_23/Y gnd 17.38fF
C85 NAND3X1_49/B gnd 49.29fF
C86 INVX1_34/A vdd 2.15fF
C87 A<2> gnd 2.06fF
C88 NAND2X1_40/B NOR2X1_12/A 2.45fF
C89 INVX4_1/Y gnd 3.58fF
C90 AOI21X1_20/Y gnd 7.49fF
C91 INVX2_7/Y vdd 4.70fF
C92 A<7> gnd 3.47fF
C93 B<4> vdd 3.15fF
C94 A<5> gnd 72.09fF
C95 B<2> vdd 2.45fF
C96 NAND2X1_24/B gnd 4.72fF
C97 vdd NAND3X1_49/C 2.85fF
C98 NAND2X1_15/Y vdd 2.96fF
C99 A<6> gnd 2.37fF
C100 vdd gnd 30.33fF
C101 AOI21X1_76/A vdd 2.30fF
C102 A<4> gnd 2.80fF
C103 NOR2X1_25/A vdd 2.37fF
C104 AND2X2_11/Y vdd 2.04fF
C105 NOR2X1_46/B gnd 5.21fF
C106 AND2X2_14/Y vdd 2.94fF
C107 AOI21X1_4/Y vdd 4.13fF
C108 NAND3X1_6/C vdd 5.85fF
C109 OAI21X1_6/C vdd 2.07fF
C110 NOR2X1_14/B vdd 2.56fF
C111 B<7> vdd 2.19fF
C112 AND2X2_3/B AND2X2_3/A 2.27fF
C113 BUFX4_3/Y BUFX4_2/Y 2.07fF
C114 gnd NAND3X1_49/Y 2.40fF
C115 OAI21X1_68/Y vdd 3.44fF
C116 AOI21X1_72/B vdd 2.01fF
C117 INVX1_48/A vdd 2.27fF
C118 gnd AOI21X1_40/Y 10.49fF
C119 B<3> vdd 3.12fF
C120 NAND2X1_45/Y vdd 2.48fF
C121 INVX2_4/Y vdd 3.07fF
C122 NOR2X1_14/B INVX2_1/Y 2.34fF
XFILL_1_1 gnd vdd FILL
XNAND3X1_36 INVX1_12/A INVX1_22/A AOI21X1_33/B gnd NAND2X1_40/A vdd NAND3X1
XNAND3X1_24 NAND3X1_24/A NAND3X1_24/B OAI21X1_9/Y gnd INVX1_9/A vdd NAND3X1
XBUFX2_11 BUFX2_11/A gnd S<10> vdd BUFX2
XAOI21X1_33 INVX1_12/A AOI21X1_33/B INVX1_22/Y gnd OAI22X1_2/C vdd AOI21X1
XNOR2X1_12 NOR2X1_12/A NOR2X1_12/B gnd INVX1_13/A vdd NOR2X1
XNAND2X1_40 NAND2X1_40/A NAND2X1_40/B gnd NOR2X1_12/B vdd NAND2X1
XINVX1_12 INVX1_12/A gnd INVX1_12/Y vdd INVX1
XNAND3X1_49 INVX1_13/Y NAND3X1_49/B NAND3X1_49/C gnd NAND3X1_49/Y vdd NAND3X1
XAOI21X1_16 NAND2X1_21/Y NAND2X1_23/Y AOI21X1_22/A gnd gnd vdd AOI21X1
XAOI21X1_22 AOI21X1_22/A NAND2X1_23/Y NOR2X1_7/Y gnd AOI21X1_22/Y vdd AOI21X1
XNAND2X1_23 NOR2X1_7/A NOR2X1_7/B gnd NAND2X1_23/Y vdd NAND2X1
XNOR2X1_7 NOR2X1_7/A NOR2X1_7/B gnd NOR2X1_7/Y vdd NOR2X1
XNAND2X1_26 NOR2X1_7/B AND2X2_5/Y gnd NAND2X1_26/Y vdd NAND2X1
XNAND2X1_25 NOR2X1_7/A NOR2X1_8/A gnd NAND2X1_25/Y vdd NAND2X1
XNAND2X1_21 NOR2X1_8/A AND2X2_5/Y gnd NAND2X1_21/Y vdd NAND2X1
XAOI21X1_13 NAND2X1_2/Y OR2X2_1/Y AND2X2_2/Y gnd NOR2X1_7/B vdd AOI21X1
XOR2X2_1 OR2X2_1/A OR2X2_1/B gnd OR2X2_1/Y vdd OR2X2
XAND2X2_2 OR2X2_1/A OR2X2_1/B gnd AND2X2_2/Y vdd AND2X2
XNAND2X1_5 NAND3X1_3/Y NAND3X1_4/Y gnd NAND2X1_5/Y vdd NAND2X1
XNAND2X1_2 NAND2X1_2/A NAND3X1_1/Y gnd NAND2X1_2/Y vdd NAND2X1
XNAND3X1_131 INVX1_57/A NAND3X1_3/B NAND3X1_3/C gnd NAND2X1_2/A vdd NAND3X1
XNAND3X1_3 INVX1_57/Y NAND3X1_3/B NAND3X1_3/C gnd NAND3X1_3/Y vdd NAND3X1
XAOI21X1_12 NAND3X1_3/B INVX1_57/Y NOR2X1_5/Y gnd AOI21X1_12/Y vdd AOI21X1
XINVX1_57 INVX1_57/A gnd INVX1_57/Y vdd INVX1
XNAND3X1_1 INVX1_57/Y NAND2X1_1/Y OAI21X1_1/Y gnd NAND3X1_1/Y vdd NAND3X1
XNAND3X1_4 INVX1_57/A NAND2X1_1/Y OAI21X1_1/Y gnd NAND3X1_4/Y vdd NAND3X1
XOAI21X1_1 INVX4_1/Y INVX4_6/Y NOR2X1_4/A gnd OAI21X1_1/Y vdd OAI21X1
XOAI21X1_126 INVX4_1/Y INVX4_6/Y NOR2X1_5/A gnd NAND3X1_3/B vdd OAI21X1
XNAND2X1_1 NOR2X1_5/A NOR2X1_4/B gnd NAND2X1_1/Y vdd NAND2X1
XAND2X2_25 B<3> A<5> gnd NOR2X1_4/B vdd AND2X2
XNOR2X1_5 NOR2X1_5/A NOR2X1_5/B gnd NOR2X1_5/Y vdd NOR2X1
XNAND2X1_127 A<4> B<4> gnd NOR2X1_5/A vdd NAND2X1
XNAND2X1_14 B<3> A<5> gnd NOR2X1_5/B vdd NAND2X1
XAND2X2_24 A<4> B<4> gnd NOR2X1_4/A vdd AND2X2
XAOI21X1_1 AND2X2_18/Y vdd AOI22X1_1/Y gnd OR2X2_1/B vdd AOI21X1
XAND2X2_1 B<2> A<7> gnd vdd vdd AND2X2
XAOI22X1_1 B<1> A<7> B<2> A<6> gnd AOI22X1_1/Y vdd AOI22X1
XAND2X2_18 B<1> A<6> gnd AND2X2_18/Y vdd AND2X2
XNAND2X1_115 B<2> A<5> gnd INVX1_52/A vdd NAND2X1
XAOI22X1_17 B<0> A<7> B<1> A<6> gnd INVX1_53/A vdd AOI22X1
XINVX1_52 INVX1_52/A gnd INVX1_52/Y vdd INVX1
XINVX1_53 INVX1_53/A gnd INVX1_53/Y vdd INVX1
XNAND3X1_109 INVX1_52/Y INVX1_53/Y AOI22X1_19/D gnd AOI21X1_82/A vdd NAND3X1
XAOI22X1_19 B<2> A<5> INVX1_53/Y AOI22X1_19/D gnd NOR3X1_1/C vdd AOI22X1
XAND2X2_23 B<1> A<7> gnd AND2X2_23/Y vdd AND2X2
XNAND2X1_116 AND2X2_22/Y AND2X2_23/Y gnd AOI22X1_19/D vdd NAND2X1
XDFFPOSX1_4 BUFX2_1/A clk NOR2X1_24/Y gnd vdd DFFPOSX1
XBUFX2_1 BUFX2_1/A gnd S<0> vdd BUFX2
XINVX1_31 vdd gnd INVX1_31/Y vdd INVX1
XNAND2X1_76 AOI22X1_9/D NAND2X1_76/B gnd NAND2X1_76/Y vdd NAND2X1
XXNOR2X1_5 XNOR2X1_5/A INVX1_31/Y gnd XNOR2X1_5/Y vdd XNOR2X1
XINVX1_29 INVX1_29/A gnd INVX1_29/Y vdd INVX1
XNOR2X1_26 NOR2X1_26/A INVX1_29/Y gnd NOR2X1_26/Y vdd NOR2X1
XDFFPOSX1_5 BUFX2_2/A clk NOR2X1_26/Y gnd vdd DFFPOSX1
XBUFX2_2 BUFX2_2/A gnd S<1> vdd BUFX2
XFILL_2_1 gnd vdd FILL
XINVX1_22 INVX1_22/A gnd INVX1_22/Y vdd INVX1
XNAND2X1_41 AOI22X1_6/D AOI22X1_6/C gnd INVX1_14/A vdd NAND2X1
XNAND3X1_39 NAND2X1_40/A NAND2X1_40/B NOR2X1_12/A gnd AOI22X1_6/D vdd NAND3X1
XAOI21X1_19 AOI21X1_19/A INVX1_9/A INVX1_6/A gnd AOI21X1_19/Y vdd AOI21X1
XNAND2X1_28 NAND3X1_22/C NAND2X1_24/A gnd INVX1_12/A vdd NAND2X1
XNAND3X1_22 INVX1_3/Y NAND3X1_22/B NAND3X1_22/C gnd NAND2X1_24/A vdd NAND3X1
XNAND2X1_16 NAND2X1_16/A NAND2X1_16/B gnd AOI21X1_22/A vdd NAND2X1
XNAND2X1_24 NAND2X1_24/A NAND2X1_24/B gnd AOI21X1_15/C vdd NAND2X1
XNAND3X1_21 NAND2X1_23/Y NAND2X1_21/Y AOI21X1_22/A gnd NAND3X1_24/A vdd NAND3X1
XOAI21X1_23 AOI21X1_15/C NOR2X1_8/Y NAND2X1_21/Y gnd OAI21X1_23/Y vdd OAI21X1
XOAI21X1_18 NOR2X1_7/Y NOR2X1_8/Y AOI21X1_15/C gnd NAND3X1_24/B vdd OAI21X1
XAOI21X1_15 NAND2X1_26/Y NAND2X1_25/Y AOI21X1_15/C gnd AOI21X1_15/Y vdd AOI21X1
XNOR2X1_8 NOR2X1_8/A AND2X2_5/Y gnd NOR2X1_8/Y vdd NOR2X1
XNAND3X1_2 NAND2X1_4/Y OR2X2_1/Y NAND2X1_2/Y gnd NAND3X1_2/Y vdd NAND3X1
XOAI21X1_13 NOR2X1_1/Y NAND2X1_5/Y NAND2X1_4/Y gnd NOR2X1_8/A vdd OAI21X1
XOAI21X1_2 NOR2X1_1/Y AND2X2_2/Y NAND2X1_5/Y gnd OAI21X1_2/Y vdd OAI21X1
XNAND2X1_4 OR2X2_1/B OR2X2_1/A gnd NAND2X1_4/Y vdd NAND2X1
XNOR2X1_1 OR2X2_1/B OR2X2_1/A gnd NOR2X1_1/Y vdd NOR2X1
XAND2X2_5 AND2X2_5/A AND2X2_5/B gnd AND2X2_5/Y vdd AND2X2
XNAND2X1_22 AND2X2_5/A AND2X2_5/B gnd NOR2X1_7/A vdd NAND2X1
XOAI21X1_10 INVX1_57/A NOR2X1_4/Y NAND3X1_3/C gnd OAI21X1_10/Y vdd OAI21X1
XNAND2X1_126 NOR2X1_4/A NOR2X1_4/B gnd NAND3X1_3/C vdd NAND2X1
XNOR2X1_4 NOR2X1_4/A NOR2X1_4/B gnd NOR2X1_4/Y vdd NOR2X1
XNAND3X1_20 gnd NAND3X1_20/B OAI21X1_17/Y gnd AND2X2_5/B vdd NAND3X1
XOAI21X1_17 AOI22X1_3/Y NOR2X1_6/Y INVX1_5/Y gnd OAI21X1_17/Y vdd OAI21X1
XNAND2X1_125 A<3> B<5> gnd INVX1_57/A vdd NAND2X1
XINVX4_6 A<5> gnd INVX4_6/Y vdd INVX4
XOAI21X1_16 AOI22X1_3/Y NOR2X1_6/Y INVX1_5/A gnd NAND3X1_18/C vdd OAI21X1
XNAND3X1_18 INVX1_4/Y NAND3X1_18/B NAND3X1_18/C gnd AND2X2_5/A vdd NAND3X1
XINVX1_4 gnd gnd INVX1_4/Y vdd INVX1
XNOR2X1_6 NOR2X1_5/B NOR2X1_6/B gnd NOR2X1_6/Y vdd NOR2X1
XNAND2X1_20 B<4> A<6> gnd NOR2X1_6/B vdd NAND2X1
XAOI22X1_3 B<3> A<6> B<4> A<5> gnd AOI22X1_3/Y vdd AOI22X1
XINVX4_5 A<6> gnd vdd vdd INVX4
XOAI21X1_14 INVX2_7/Y vdd vdd gnd gnd vdd OAI21X1
XOAI22X1_1 OAI22X1_1/A NAND2X1_3/Y INVX1_52/A INVX1_53/A gnd OR2X2_1/A vdd OAI22X1
XNAND2X1_3 B<1> A<7> gnd NAND2X1_3/Y vdd NAND2X1
XNAND2X1_117 B<1> A<6> gnd NAND3X1_110/C vdd NAND2X1
XNAND3X1_110 B<0> A<7> NAND3X1_110/C gnd AOI21X1_70/A vdd NAND3X1
XAOI21X1_70 AOI21X1_70/A AOI21X1_70/B INVX1_52/A gnd NOR3X1_1/B vdd AOI21X1
XNAND3X1_112 INVX1_52/A AOI21X1_70/A AOI21X1_70/B gnd AOI21X1_82/B vdd NAND3X1
XNAND3X1_111 B<1> A<6> NAND2X1_118/Y gnd AOI21X1_70/B vdd NAND3X1
XNAND2X1_118 B<0> A<7> gnd NAND2X1_118/Y vdd NAND2X1
XNAND3X1_91 B<1> A<5> OAI22X1_1/A gnd NAND3X1_91/Y vdd NAND3X1
XNAND2X1_105 B<0> A<6> gnd OAI22X1_1/A vdd NAND2X1
XAND2X2_22 B<0> A<6> gnd AND2X2_22/Y vdd AND2X2
XINVX4_1 B<3> gnd INVX4_1/Y vdd INVX4
XNOR2X1_24 gnd INVX2_4/Y gnd NOR2X1_24/Y vdd NOR2X1
XINVX2_4 B<0> gnd INVX2_4/Y vdd INVX2
XINVX2_7 B<1> gnd INVX2_7/Y vdd INVX2
XNOR2X1_28 gnd INVX2_7/Y gnd NOR2X1_25/B vdd NOR2X1
XNOR2X1_25 NOR2X1_25/A NOR2X1_25/B gnd NOR2X1_26/A vdd NOR2X1
XNAND2X1_72 NOR2X1_25/A NOR2X1_25/B gnd INVX1_29/A vdd NAND2X1
XNAND2X1_74 INVX1_32/Y NOR2X1_25/A gnd NAND2X1_76/B vdd NAND2X1
XNOR2X1_30 INVX1_29/A XNOR2X1_5/Y gnd INVX1_33/A vdd NOR2X1
XXNOR2X1_4 XNOR2X1_5/Y INVX1_29/Y gnd XNOR2X1_4/Y vdd XNOR2X1
XDFFPOSX1_6 BUFX2_3/A clk XNOR2X1_4/Y gnd vdd DFFPOSX1
XBUFX2_3 BUFX2_3/A gnd S<2> vdd BUFX2
XFILL_3_4 gnd vdd FILL
XFILL_3_3 gnd vdd FILL
XFILL_3_2 gnd vdd FILL
XFILL_3_1 gnd vdd FILL
XNAND3X1_15 vdd NAND3X1_22/B NAND3X1_22/C gnd NAND2X1_16/A vdd NAND3X1
XINVX1_3 vdd gnd INVX1_3/Y vdd INVX1
XNAND3X1_16 INVX1_3/Y NAND2X1_15/Y OAI21X1_12/Y gnd NAND2X1_16/B vdd NAND3X1
XNAND3X1_23 vdd NAND2X1_15/Y OAI21X1_12/Y gnd NAND2X1_24/B vdd NAND3X1
XNOR2X1_9 NOR2X1_9/A NOR2X1_9/B gnd NOR2X1_9/Y vdd NOR2X1
XNAND2X1_9 NOR2X1_9/A NOR2X1_9/B gnd NAND2X1_9/Y vdd NAND2X1
XNAND2X1_6 OAI21X1_2/Y NAND3X1_2/Y gnd NOR2X1_9/B vdd NAND2X1
XAOI21X1_11 NAND3X1_2/Y OAI21X1_2/Y NAND3X1_6/C gnd OAI21X1_9/A vdd AOI21X1
XNAND2X1_7 NAND3X1_6/C NOR2X1_9/B gnd NAND2X1_7/Y vdd NAND2X1
XNAND3X1_5 NAND3X1_2/Y OAI21X1_2/Y NOR2X1_9/A gnd NAND3X1_5/Y vdd NAND3X1
XNAND3X1_6 NAND3X1_2/Y OAI21X1_2/Y NAND3X1_6/C gnd NAND3X1_6/Y vdd NAND3X1
XNAND2X1_35 NAND2X1_34/Y AND2X2_5/A gnd OR2X2_2/A vdd NAND2X1
XNAND2X1_13 NOR2X1_3/Y OAI21X1_10/Y gnd NAND3X1_22/C vdd NAND2X1
XNAND2X1_15 NOR2X1_3/Y AOI21X1_12/Y gnd NAND2X1_15/Y vdd NAND2X1
XNOR2X1_3 vdd BUFX4_1/Y gnd NOR2X1_3/Y vdd NOR2X1
XOAI21X1_12 vdd BUFX4_3/Y OAI21X1_10/Y gnd OAI21X1_12/Y vdd OAI21X1
XOAI21X1_11 vdd BUFX4_2/Y AOI21X1_12/Y gnd NAND3X1_22/B vdd OAI21X1
XAOI22X1_5 NOR2X1_4/B gnd INVX1_5/Y AOI22X1_5/D gnd AOI22X1_5/Y vdd AOI22X1
XNAND2X1_18 NOR2X1_4/B gnd gnd NAND3X1_19/C vdd NAND2X1
XNAND3X1_17 INVX1_5/Y AOI22X1_5/D NAND3X1_19/C gnd NAND3X1_18/B vdd NAND3X1
XNAND3X1_19 INVX1_5/A AOI22X1_5/D NAND3X1_19/C gnd NAND3X1_20/B vdd NAND3X1
XOAI21X1_24 INVX1_5/A AOI22X1_3/Y OAI21X1_24/C gnd OAI21X1_24/Y vdd OAI21X1
XINVX1_5 INVX1_5/A gnd INVX1_5/Y vdd INVX1
XNAND2X1_36 B<4> A<7> gnd NOR2X1_14/B vdd NAND2X1
XNAND2X1_12 A<2> B<7> gnd vdd vdd NAND2X1
XAND2X2_4 B<4> A<6> gnd gnd vdd AND2X2
XNAND2X1_17 A<4> B<5> gnd INVX1_5/A vdd NAND2X1
XAND2X2_20 B<3> A<4> gnd AND2X2_20/Y vdd AND2X2
XNAND2X1_34 AND2X2_18/Y vdd gnd NAND2X1_34/Y vdd NAND2X1
XOAI21X1_125 OAI21X1_125/A AOI21X1_82/Y AOI21X1_72/B gnd NAND3X1_6/C vdd OAI21X1
XNAND3X1_114 AOI21X1_2/A AOI21X1_72/B AOI21X1_2/B gnd AOI21X1_81/A vdd NAND3X1
XAOI21X1_2 AOI21X1_2/A AOI21X1_2/B NOR3X1_1/Y gnd NOR2X1_9/A vdd AOI21X1
XAOI21X1_72 AOI21X1_2/B AOI21X1_72/B AOI21X1_2/A gnd NOR3X1_2/B vdd AOI21X1
XNOR3X1_1 NOR3X1_1/A NOR3X1_1/B NOR3X1_1/C gnd NOR3X1_1/Y vdd NOR3X1
XOAI21X1_110 NOR3X1_1/B NOR3X1_1/C NOR3X1_1/A gnd AOI21X1_2/B vdd OAI21X1
XOAI21X1_111 NOR3X1_1/B NOR3X1_1/C AOI21X1_82/C gnd AOI22X1_20/D vdd OAI21X1
XAOI21X1_82 AOI21X1_82/A AOI21X1_82/B AOI21X1_82/C gnd AOI21X1_82/Y vdd AOI21X1
XNAND3X1_113 AOI21X1_82/B AOI21X1_82/A AOI21X1_82/C gnd AOI21X1_72/B vdd NAND3X1
XNAND3X1_117 AOI21X1_82/B NOR3X1_1/A AOI21X1_82/A gnd AOI22X1_20/C vdd NAND3X1
XOAI21X1_109 INVX1_44/A AND2X2_21/Y AOI22X1_14/D gnd AOI21X1_82/C vdd OAI21X1
XNAND2X1_103 AND2X2_14/Y AND2X2_18/Y gnd AOI22X1_14/D vdd NAND2X1
XAND2X2_21 INVX1_45/A OAI22X1_1/A gnd AND2X2_21/Y vdd AND2X2
XNAND2X1_104 B<1> A<5> gnd INVX1_45/A vdd NAND2X1
XNAND2X1_96 B<0> A<5> gnd NAND2X1_96/Y vdd NAND2X1
XAND2X2_14 B<0> A<5> gnd AND2X2_14/Y vdd AND2X2
XAND2X2_13 A<4> B<1> gnd AND2X2_13/Y vdd AND2X2
XINVX4_2 A<3> gnd vdd vdd INVX4
XNOR2X1_29 gnd INVX1_30/Y gnd vdd vdd NOR2X1
XINVX1_30 B<2> gnd INVX1_30/Y vdd INVX1
XNOR2X1_27 INVX2_4/Y vdd gnd NOR2X1_25/A vdd NOR2X1
XOAI21X1_60 INVX2_7/Y vdd OAI22X1_5/A gnd AOI22X1_9/D vdd OAI21X1
XAOI22X1_9 NOR2X1_25/A INVX1_32/Y vdd AOI22X1_9/D gnd INVX1_34/A vdd AOI22X1
XINVX1_32 AND2X2_9/A gnd INVX1_32/Y vdd INVX1
XNAND2X1_75 B<0> A<2> gnd OAI22X1_5/A vdd NAND2X1
XNAND2X1_83 B<0> A<3> gnd AND2X2_9/B vdd NAND2X1
XAND2X2_9 AND2X2_9/A AND2X2_9/B gnd AND2X2_9/Y vdd AND2X2
XNOR2X1_36 AND2X2_9/A AND2X2_9/B gnd NOR2X1_36/Y vdd NOR2X1
XNAND2X1_73 B<1> A<2> gnd AND2X2_9/A vdd NAND2X1
XFILL_4_2 gnd vdd FILL
XFILL_4_1 gnd vdd FILL
XOAI21X1_19 gnd AOI21X1_15/Y AOI21X1_14/Y gnd AOI21X1_19/A vdd OAI21X1
XOAI21X1_20 gnd AOI21X1_15/Y OAI21X1_9/Y gnd OAI21X1_20/Y vdd OAI21X1
XAOI21X1_14 NAND2X1_8/Y NAND2X1_9/Y NOR2X1_9/Y gnd AOI21X1_14/Y vdd AOI21X1
XNAND3X1_7 NAND2X1_8/Y NAND3X1_6/Y NAND2X1_9/Y gnd NAND3X1_7/Y vdd NAND3X1
XOAI21X1_9 OAI21X1_9/A AND2X2_3/Y NAND3X1_6/Y gnd OAI21X1_9/Y vdd OAI21X1
XAND2X2_3 AND2X2_3/A AND2X2_3/B gnd AND2X2_3/Y vdd AND2X2
XNAND2X1_8 AND2X2_3/B AND2X2_3/A gnd NAND2X1_8/Y vdd NAND2X1
XNAND3X1_8 AND2X2_3/Y NAND2X1_7/Y NAND3X1_5/Y gnd NAND3X1_8/Y vdd NAND3X1
XAOI22X1_2 AND2X2_3/B AND2X2_3/A NAND2X1_7/Y NAND3X1_5/Y gnd AOI22X1_2/Y vdd AOI22X1
XNAND3X1_31 NAND2X1_34/Y AND2X2_5/A OR2X2_2/B gnd gnd vdd NAND3X1
XXOR2X1_2 XOR2X1_2/A XOR2X1_2/B gnd OR2X2_2/B vdd XOR2X1
XOAI21X1_25 INVX4_3/Y BUFX4_1/Y AOI22X1_5/Y gnd OAI21X1_25/Y vdd OAI21X1
XNOR2X1_11 INVX4_6/Y INVX2_1/Y gnd XOR2X1_2/B vdd NOR2X1
XAOI21X1_27 OAI21X1_26/Y XOR2X1_2/B NOR2X1_14/Y gnd INVX1_18/A vdd AOI21X1
XOAI21X1_27 NOR2X1_14/A NOR2X1_14/B OAI21X1_26/Y gnd XOR2X1_2/A vdd OAI21X1
XNOR2X1_14 NOR2X1_14/A NOR2X1_14/B gnd NOR2X1_14/Y vdd NOR2X1
XOAI21X1_15 INVX2_9/Y INVX4_6/Y NOR2X1_14/A gnd AOI22X1_5/D vdd OAI21X1
XNAND2X1_30 NOR2X1_10/Y OAI21X1_24/Y gnd NAND2X1_30/Y vdd NAND2X1
XNOR2X1_10 INVX4_3/Y BUFX4_4/Y gnd NOR2X1_10/Y vdd NOR2X1
XOAI21X1_26 INVX4_1/Y INVX2_2/Y OAI21X1_26/C gnd OAI21X1_26/Y vdd OAI21X1
XINVX2_2 A<7> gnd INVX2_2/Y vdd INVX2
XINVX2_1 B<5> gnd INVX2_1/Y vdd INVX2
XOAI22X1_6 INVX4_1/Y INVX4_3/Y vdd INVX2_9/Y gnd OAI22X1_6/Y vdd OAI22X1
XNAND2X1_19 B<3> A<6> gnd NOR2X1_14/A vdd NAND2X1
XAOI22X1_22 AND2X2_16/Y NOR2X1_4/A INVX1_51/Y OAI22X1_6/Y gnd AOI22X1_22/Y vdd AOI22X1
XINVX1_51 INVX1_51/A gnd INVX1_51/Y vdd INVX1
XNAND3X1_115 INVX1_51/Y OAI22X1_6/Y NAND3X1_107/C gnd NAND2X1_119/A vdd NAND3X1
XNAND3X1_107 INVX1_51/A OAI22X1_6/Y NAND3X1_107/C gnd AOI22X1_20/A vdd NAND3X1
XNAND2X1_119 NAND2X1_119/A NAND3X1_116/Y gnd OAI21X1_125/A vdd NAND2X1
XNAND3X1_116 INVX1_51/A OAI21X1_107/Y NAND3X1_108/C gnd NAND3X1_116/Y vdd NAND3X1
XNAND3X1_108 INVX1_51/Y OAI21X1_107/Y NAND3X1_108/C gnd AOI22X1_20/B vdd NAND3X1
XOAI21X1_107 vdd INVX2_9/Y AND2X2_20/Y gnd OAI21X1_107/Y vdd OAI21X1
XNAND2X1_114 AOI22X1_20/A AOI22X1_20/B gnd AOI21X1_2/A vdd NAND2X1
XAOI22X1_20 AOI22X1_20/A AOI22X1_20/B AOI22X1_20/C AOI22X1_20/D gnd NOR3X1_2/A vdd
+ AOI22X1
XNAND3X1_118 OAI21X1_125/A AOI22X1_20/C AOI22X1_20/D gnd AOI21X1_81/B vdd NAND3X1
XNAND2X1_102 A<4> B<2> gnd INVX1_44/A vdd NAND2X1
XNAND3X1_90 B<0> A<6> INVX1_45/A gnd NAND3X1_90/Y vdd NAND3X1
XINVX1_44 INVX1_44/A gnd INVX1_44/Y vdd INVX1
XNAND3X1_89 INVX1_44/Y gnd AOI22X1_14/D gnd NAND3X1_89/Y vdd NAND3X1
XAOI22X1_18 AND2X2_14/Y AND2X2_18/Y INVX1_44/Y gnd gnd NOR3X1_1/A vdd AOI22X1
XAOI22X1_14 A<4> B<2> gnd AOI22X1_14/D gnd NOR3X1_9/C vdd AOI22X1
XOAI21X1_94 INVX2_4/Y vdd INVX1_45/A gnd gnd vdd OAI21X1
XAOI22X1_12 A<4> B<1> B<0> A<5> gnd AOI22X1_12/Y vdd AOI22X1
XAND2X2_11 A<4> B<0> gnd AND2X2_11/Y vdd AND2X2
XINVX4_3 A<4> gnd INVX4_3/Y vdd INVX4
XNAND2X1_86 A<4> B<0> gnd NOR2X1_35/B vdd NAND2X1
XAND2X2_10 B<1> A<3> gnd AND2X2_10/Y vdd AND2X2
XOAI21X1_71 INVX4_3/Y INVX2_4/Y AND2X2_10/Y gnd OAI21X1_71/Y vdd OAI21X1
XOAI21X1_68 INVX4_3/Y INVX2_4/Y OAI22X1_5/B gnd OAI21X1_68/Y vdd OAI21X1
XOAI21X1_61 INVX2_4/Y vdd AND2X2_9/A gnd AOI21X1_44/A vdd OAI21X1
XNAND2X1_78 B<1> A<3> gnd OAI22X1_5/B vdd NAND2X1
XOAI22X1_5 OAI22X1_5/A OAI22X1_5/B INVX1_35/A AND2X2_9/Y gnd OAI22X1_5/Y vdd OAI22X1
XOAI21X1_62 OAI22X1_5/A OAI22X1_5/B AOI21X1_44/A gnd XNOR2X1_6/A vdd OAI21X1
XAOI21X1_44 AOI21X1_44/A INVX1_35/Y NOR2X1_36/Y gnd NOR3X1_5/A vdd AOI21X1
XINVX1_35 INVX1_35/A gnd INVX1_35/Y vdd INVX1
XFILL_5_2 gnd vdd FILL
XFILL_5_1 gnd vdd FILL
XAOI21X1_18 NAND3X1_27/C OAI21X1_20/Y INVX1_6/Y gnd AOI21X1_18/Y vdd AOI21X1
XNAND3X1_27 INVX1_6/Y OAI21X1_20/Y NAND3X1_27/C gnd NAND3X1_27/Y vdd NAND3X1
XOAI21X1_29 AOI21X1_24/Y OAI21X1_30/B AOI21X1_22/Y gnd AOI21X1_33/B vdd OAI21X1
XOAI21X1_30 AOI21X1_24/Y OAI21X1_30/B OAI21X1_23/Y gnd OAI21X1_30/Y vdd OAI21X1
XAOI21X1_24 INVX1_16/A gnd NAND2X1_33/Y gnd AOI21X1_24/Y vdd AOI21X1
XAOI21X1_3 NAND2X1_9/Y NAND3X1_6/Y NAND2X1_8/Y gnd AOI21X1_3/Y vdd AOI21X1
XINVX1_21 gnd gnd INVX1_21/Y vdd INVX1
XNAND2X1_37 OR2X2_2/A INVX1_11/Y gnd INVX1_16/A vdd NAND2X1
XINVX1_11 OR2X2_2/B gnd INVX1_11/Y vdd INVX1
XNAND2X1_39 OR2X2_2/B OR2X2_2/A gnd NAND2X1_39/Y vdd NAND2X1
XOR2X2_2 OR2X2_2/A OR2X2_2/B gnd OR2X2_2/Y vdd OR2X2
XNAND2X1_33 NAND3X1_30/Y NAND2X1_32/Y gnd NAND2X1_33/Y vdd NAND2X1
XNAND2X1_32 INVX1_10/Y NAND2X1_31/Y gnd NAND2X1_32/Y vdd NAND2X1
XINVX1_10 INVX1_10/A gnd INVX1_10/Y vdd INVX1
XNAND3X1_33 INVX1_10/Y NAND2X1_30/Y OAI21X1_25/Y gnd NAND3X1_33/Y vdd NAND3X1
XNAND3X1_30 INVX1_10/A NAND2X1_30/Y OAI21X1_25/Y gnd NAND3X1_30/Y vdd NAND3X1
XNAND2X1_31 NAND2X1_30/Y OAI21X1_25/Y gnd NAND2X1_31/Y vdd NAND2X1
XOAI21X1_37 INVX2_1/Y vdd NOR2X1_14/B gnd OAI21X1_37/Y vdd OAI21X1
XNAND2X1_29 A<3> B<7> gnd INVX1_10/A vdd NAND2X1
XOAI21X1_8 INVX1_56/A OAI21X1_8/B OAI21X1_8/C gnd INVX1_6/A vdd OAI21X1
XNAND2X1_11 NAND2X1_11/A OAI21X1_8/C gnd OAI21X1_8/B vdd NAND2X1
XNAND3X1_129 INVX1_56/A NAND2X1_11/A OAI21X1_8/C gnd AND2X2_3/B vdd NAND3X1
XNAND3X1_130 INVX1_56/Y NAND2X1_124/Y OAI21X1_124/Y gnd AND2X2_3/A vdd NAND3X1
XINVX1_56 INVX1_56/A gnd INVX1_56/Y vdd INVX1
XNAND2X1_123 NOR2X1_47/Y OAI21X1_122/Y gnd OAI21X1_8/C vdd NAND2X1
XNAND2X1_124 NOR2X1_47/Y AOI22X1_22/Y gnd NAND2X1_124/Y vdd NAND2X1
XNOR2X1_47 INVX4_4/Y BUFX4_2/Y gnd NOR2X1_47/Y vdd NOR2X1
XOAI21X1_123 INVX4_4/Y BUFX4_3/Y AOI22X1_22/Y gnd NAND2X1_11/A vdd OAI21X1
XOAI21X1_124 INVX4_4/Y BUFX4_4/Y OAI21X1_122/Y gnd OAI21X1_124/Y vdd OAI21X1
XOAI21X1_122 INVX1_51/A NOR2X1_48/Y NAND3X1_107/C gnd OAI21X1_122/Y vdd OAI21X1
XNOR2X1_48 AND2X2_19/Y AND2X2_20/Y gnd NOR2X1_48/Y vdd NOR2X1
XNAND2X1_113 AND2X2_19/Y AND2X2_20/Y gnd NAND3X1_107/C vdd NAND2X1
XAND2X2_16 B<3> A<3> gnd AND2X2_16/Y vdd AND2X2
XOAI21X1_108 INVX4_1/Y INVX4_3/Y AND2X2_19/Y gnd NAND3X1_108/C vdd OAI21X1
XAND2X2_19 A<3> B<4> gnd AND2X2_19/Y vdd AND2X2
XNOR3X1_2 NOR3X1_2/A NOR3X1_2/B NOR3X1_2/C gnd vdd vdd NOR3X1
XINVX4_4 A<2> gnd INVX4_4/Y vdd INVX4
XNAND3X1_92 INVX1_44/A NAND3X1_90/Y NAND3X1_91/Y gnd NAND3X1_95/A vdd NAND3X1
XAOI21X1_61 NAND3X1_90/Y NAND3X1_91/Y INVX1_44/A gnd NOR3X1_9/B vdd AOI21X1
XNOR3X1_9 NOR3X1_9/A NOR3X1_9/B NOR3X1_9/C gnd NOR3X1_9/Y vdd NOR3X1
XINVX1_45 INVX1_45/A gnd INVX1_45/Y vdd INVX1
XAOI22X1_13 AND2X2_11/Y INVX1_45/Y INVX1_42/Y AOI22X1_10/C gnd NOR3X1_9/A vdd AOI22X1
XOAI21X1_79 INVX4_3/Y INVX2_7/Y NAND2X1_96/Y gnd AOI22X1_10/C vdd OAI21X1
XNAND2X1_95 AND2X2_13/Y AND2X2_14/Y gnd AOI22X1_10/D vdd NAND2X1
XNAND2X1_97 NAND2X1_96/Y AND2X2_13/Y gnd NAND2X1_97/Y vdd NAND2X1
XOAI21X1_80 INVX4_3/Y INVX2_7/Y AND2X2_14/Y gnd OAI21X1_80/Y vdd OAI21X1
XNAND2X1_94 A<3> B<2> gnd INVX1_42/A vdd NAND2X1
XAOI22X1_10 A<3> B<2> AOI22X1_10/C AOI22X1_10/D gnd NOR3X1_7/B vdd AOI22X1
XNAND2X1_85 AND2X2_10/Y AND2X2_11/Y gnd NAND2X1_85/Y vdd NAND2X1
XOAI21X1_70 INVX2_7/Y vdd AND2X2_11/Y gnd AOI21X1_45/A vdd OAI21X1
XINVX2_5 A<1> gnd vdd vdd INVX2
XAND2X2_12 OAI22X1_5/B NOR2X1_35/B gnd AND2X2_12/Y vdd AND2X2
XNOR2X1_35 OAI22X1_5/B NOR2X1_35/B gnd NOR2X1_35/Y vdd NOR2X1
XAOI21X1_45 AOI21X1_45/A OAI21X1_71/Y INVX1_36/A gnd NOR3X1_5/C vdd AOI21X1
XNAND2X1_84 B<2> A<2> gnd INVX1_36/A vdd NAND2X1
XNAND2X1_77 B<2> A<1> gnd INVX1_35/A vdd NAND2X1
XXNOR2X1_6 XNOR2X1_6/A INVX1_35/Y gnd XNOR2X1_6/Y vdd XNOR2X1
XNAND3X1_38 INVX1_12/Y NAND3X1_37/Y OAI21X1_30/Y gnd NAND2X1_40/B vdd NAND3X1
XOAI21X1_33 INVX1_12/Y AOI21X1_26/Y INVX1_22/A gnd OAI21X1_33/Y vdd OAI21X1
XNAND3X1_37 NAND3X1_32/Y AOI21X1_22/Y NAND3X1_34/Y gnd NAND3X1_37/Y vdd NAND3X1
XNAND3X1_35 NAND3X1_32/Y NAND3X1_34/Y OAI21X1_23/Y gnd INVX1_22/A vdd NAND3X1
XAOI21X1_26 NAND3X1_34/Y NAND3X1_32/Y OAI21X1_23/Y gnd AOI21X1_26/Y vdd AOI21X1
XNAND3X1_32 INVX1_16/A gnd NAND2X1_33/Y gnd NAND3X1_32/Y vdd NAND3X1
XINVX1_16 INVX1_16/A gnd INVX1_16/Y vdd INVX1
XOAI21X1_40 INVX1_21/Y NAND2X1_38/Y INVX1_16/A gnd OAI21X1_40/Y vdd OAI21X1
XAOI21X1_23 OR2X2_2/Y NAND2X1_39/Y NAND2X1_38/Y gnd OAI21X1_30/B vdd AOI21X1
XNAND3X1_34 NAND2X1_39/Y OR2X2_2/Y NAND2X1_38/Y gnd NAND3X1_34/Y vdd NAND3X1
XNAND3X1_9 NAND3X1_7/Y NAND3X1_8/Y AOI21X1_4/Y gnd NAND3X1_9/Y vdd NAND3X1
XOAI21X1_34 INVX1_10/A NAND2X1_31/Y NAND2X1_30/Y gnd INVX1_15/A vdd OAI21X1
XNAND2X1_38 NAND3X1_33/Y OAI21X1_28/Y gnd NAND2X1_38/Y vdd NAND2X1
XOAI21X1_28 vdd INVX2_3/Y NAND2X1_31/Y gnd OAI21X1_28/Y vdd OAI21X1
XNOR2X1_13 INVX4_3/Y INVX2_3/Y gnd INVX1_17/A vdd NOR2X1
XOAI21X1_36 INVX4_6/Y BUFX4_3/Y INVX1_18/A gnd vdd vdd OAI21X1
XNAND2X1_46 OAI21X1_37/Y NAND2X1_45/Y gnd INVX1_20/A vdd NAND2X1
XOAI21X1_35 INVX4_6/Y BUFX4_2/Y INVX1_18/Y gnd OAI21X1_35/Y vdd OAI21X1
XINVX1_18 INVX1_18/A gnd INVX1_18/Y vdd INVX1
XINVX2_3 B<7> gnd INVX2_3/Y vdd INVX2
XOAI21X1_47 INVX4_6/Y INVX2_3/Y OR2X2_3/A gnd NAND3X1_50/B vdd OAI21X1
XOAI21X1_48 INVX2_1/Y INVX2_2/Y NAND2X1_52/Y gnd OAI21X1_48/Y vdd OAI21X1
XNAND2X1_52 NAND3X1_50/B OR2X2_3/Y gnd NAND2X1_52/Y vdd NAND2X1
XNOR2X1_15 INVX2_1/Y INVX2_2/Y gnd NOR2X1_15/Y vdd NOR2X1
XNAND3X1_50 NOR2X1_15/Y NAND3X1_50/B OR2X2_3/Y gnd OR2X2_6/A vdd NAND3X1
XNAND2X1_45 gnd NOR2X1_15/Y gnd NAND2X1_45/Y vdd NAND2X1
XINVX2_9 B<4> gnd INVX2_9/Y vdd INVX2
XNAND2X1_122 A<1> B<7> gnd INVX1_56/A vdd NAND2X1
XNAND2X1_112 A<2> B<5> gnd INVX1_51/A vdd NAND2X1
XAOI21X1_4 AOI21X1_4/A AOI21X1_4/B vdd gnd AOI21X1_4/Y vdd AOI21X1
XAOI21X1_81 AOI21X1_81/A AOI21X1_81/B AOI21X1_81/C gnd AOI21X1_81/Y vdd AOI21X1
XNAND3X1_119 AOI21X1_81/A AOI21X1_81/B AOI21X1_81/C gnd AOI21X1_75/B vdd NAND3X1
XNAND3X1_122 AOI21X1_81/A AOI21X1_81/B NOR3X1_2/C gnd AOI21X1_74/B vdd NAND3X1
XOAI21X1_114 NOR3X1_2/A NOR3X1_2/B AOI21X1_81/C gnd AOI21X1_74/A vdd OAI21X1
XOAI21X1_112 NOR3X1_2/A NOR3X1_2/B NOR3X1_2/C gnd AOI21X1_4/B vdd OAI21X1
XOAI21X1_106 NAND3X1_96/A AOI21X1_69/Y NAND3X1_93/Y gnd AOI21X1_81/C vdd OAI21X1
XAOI21X1_69 NAND3X1_89/Y NAND3X1_95/A OAI21X1_93/Y gnd AOI21X1_69/Y vdd AOI21X1
XNAND3X1_93 NAND3X1_95/A OAI21X1_93/Y NAND3X1_89/Y gnd NAND3X1_93/Y vdd NAND3X1
XAOI21X1_71 AND2X2_17/Y OAI21X1_95/Y NOR3X1_9/Y gnd NOR3X1_2/C vdd AOI21X1
XNAND3X1_95 NAND3X1_95/A NOR3X1_9/A NAND3X1_89/Y gnd NAND3X1_95/Y vdd NAND3X1
XOAI21X1_95 NOR3X1_9/B NOR3X1_9/C NOR3X1_9/A gnd OAI21X1_95/Y vdd OAI21X1
XOAI21X1_96 NOR3X1_9/B NOR3X1_9/C OAI21X1_93/Y gnd OAI21X1_96/Y vdd OAI21X1
XOAI21X1_93 INVX1_42/A AOI22X1_12/Y AOI22X1_10/D gnd OAI21X1_93/Y vdd OAI21X1
XINVX1_42 INVX1_42/A gnd INVX1_42/Y vdd INVX1
XNAND3X1_67 INVX1_42/Y AOI22X1_10/C AOI22X1_10/D gnd NAND3X1_67/Y vdd NAND3X1
XAOI21X1_53 OAI21X1_80/Y NAND2X1_97/Y INVX1_42/A gnd AOI21X1_53/Y vdd AOI21X1
XNAND3X1_68 INVX1_42/A NAND2X1_97/Y OAI21X1_80/Y gnd vdd vdd NAND3X1
XOAI21X1_78 INVX1_36/A AND2X2_12/Y NAND2X1_85/Y gnd vdd vdd OAI21X1
XOAI21X1_69 NOR2X1_35/Y AND2X2_12/Y INVX1_36/A gnd OAI21X1_69/Y vdd OAI21X1
XAOI21X1_52 OAI21X1_68/Y INVX1_36/Y NOR2X1_35/Y gnd NOR3X1_7/A vdd AOI21X1
XNAND3X1_61 INVX1_36/Y OAI21X1_68/Y NAND2X1_85/Y gnd NAND3X1_61/Y vdd NAND3X1
XAOI21X1_46 NAND2X1_85/Y OAI21X1_68/Y INVX1_36/Y gnd NOR3X1_5/B vdd AOI21X1
XINVX1_36 INVX1_36/A gnd INVX1_36/Y vdd INVX1
XOAI21X1_72 NOR3X1_5/B NOR3X1_5/C NOR3X1_5/A gnd OAI21X1_72/Y vdd OAI21X1
XNOR3X1_5 NOR3X1_5/A NOR3X1_5/B NOR3X1_5/C gnd NOR3X1_5/Y vdd NOR3X1
XXNOR2X1_7 XNOR2X1_6/A INVX1_35/A gnd XNOR2X1_7/Y vdd XNOR2X1
XAOI21X1_25 INVX1_6/A AOI21X1_19/A INVX1_9/Y gnd NOR2X1_12/A vdd AOI21X1
XINVX1_9 INVX1_9/A gnd INVX1_9/Y vdd INVX1
XNAND3X1_25 INVX1_6/A INVX1_9/A AOI21X1_19/A gnd NAND3X1_25/Y vdd NAND3X1
XOAI21X1_41 AOI21X1_32/Y OAI21X1_41/B OAI21X1_33/Y gnd AOI22X1_6/A vdd OAI21X1
XAOI21X1_32 NAND3X1_45/C NAND3X1_44/Y INVX1_15/A gnd AOI21X1_32/Y vdd AOI21X1
XNAND3X1_45 INVX1_15/A NAND3X1_44/Y NAND3X1_45/C gnd OAI21X1_43/C vdd NAND3X1
XOAI21X1_39 INVX1_16/Y OAI21X1_30/B NAND2X1_47/Y gnd OAI21X1_39/Y vdd OAI21X1
XAOI21X1_30 NAND2X1_33/Y gnd INVX1_16/Y gnd AOI21X1_30/Y vdd AOI21X1
XNAND3X1_44 OAI21X1_38/Y OR2X2_4/B OAI21X1_40/Y gnd NAND3X1_44/Y vdd NAND3X1
XNAND2X1_47 OR2X2_4/B OAI21X1_38/Y gnd NAND2X1_47/Y vdd NAND2X1
XAOI21X1_10 NAND3X1_8/Y NAND3X1_7/Y OAI21X1_3/C gnd OAI21X1_7/B vdd AOI21X1
XNAND3X1_10 NAND3X1_7/Y NAND3X1_8/Y OAI21X1_3/C gnd INVX1_8/A vdd NAND3X1
XOAI21X1_3 AOI21X1_3/Y AOI22X1_2/Y OAI21X1_3/C gnd OAI21X1_3/Y vdd OAI21X1
XOAI21X1_4 AOI22X1_2/Y AOI21X1_3/Y AOI21X1_4/Y gnd OAI21X1_4/Y vdd OAI21X1
XOAI21X1_38 OAI21X1_38/A AOI21X1_28/Y OAI21X1_38/C gnd OAI21X1_38/Y vdd OAI21X1
XINVX1_17 INVX1_17/A gnd INVX1_17/Y vdd INVX1
XAOI21X1_28 OAI21X1_35/Y NAND2X1_43/Y INVX1_17/Y gnd AOI21X1_28/Y vdd AOI21X1
XNAND3X1_41 INVX1_17/Y NAND2X1_43/Y OAI21X1_35/Y gnd NAND3X1_41/Y vdd NAND3X1
XNAND2X1_43 INVX1_19/Y INVX1_18/A gnd NAND2X1_43/Y vdd NAND2X1
XNAND2X1_44 INVX1_19/Y INVX1_18/Y gnd NAND2X1_44/Y vdd NAND2X1
XINVX1_19 INVX1_19/A gnd INVX1_19/Y vdd INVX1
XOAI21X1_45 vdd BUFX4_4/Y NAND2X1_45/Y gnd OAI21X1_46/C vdd OAI21X1
XOAI21X1_46 BUFX4_1/Y NAND2X1_45/Y OAI21X1_46/C gnd OR2X2_3/A vdd OAI21X1
XOR2X2_3 OR2X2_3/A OR2X2_3/B gnd OR2X2_3/Y vdd OR2X2
XNAND2X1_51 A<5> B<7> gnd OR2X2_3/B vdd NAND2X1
XOAI21X1_54 BUFX4_2/Y NAND2X1_45/Y OR2X2_3/Y gnd XOR2X1_3/B vdd OAI21X1
XNAND2X1_109 A<0> B<7> gnd gnd vdd NAND2X1
XOAI21X1_121 AOI21X1_74/C AOI21X1_81/Y AOI21X1_75/B gnd OAI21X1_3/C vdd OAI21X1
XNAND2X1_89 A<0> B<5> gnd INVX1_41/A vdd NAND2X1
XNAND2X1_100 A<1> B<5> gnd INVX1_43/A vdd NAND2X1
XAND2X2_15 A<2> B<4> gnd NOR2X1_43/A vdd AND2X2
XNOR2X1_43 NOR2X1_43/A AND2X2_16/Y gnd NOR2X1_43/Y vdd NOR2X1
XNAND2X1_101 NOR2X1_43/A AND2X2_16/Y gnd NAND3X1_87/C vdd NAND2X1
XOAI21X1_91 INVX4_4/Y INVX2_9/Y OAI21X1_91/C gnd vdd vdd OAI21X1
XOAI21X1_92 INVX4_1/Y vdd NOR2X1_43/A gnd NAND3X1_88/C vdd OAI21X1
XNAND3X1_88 INVX1_43/A vdd NAND3X1_88/C gnd AND2X2_17/A vdd NAND3X1
XNAND2X1_106 AND2X2_17/B AND2X2_17/A gnd NAND3X1_96/A vdd NAND2X1
XAND2X2_17 AND2X2_17/A AND2X2_17/B gnd AND2X2_17/Y vdd AND2X2
XNAND3X1_94 NAND3X1_93/Y AND2X2_17/Y OAI21X1_95/Y gnd NAND3X1_94/Y vdd NAND3X1
XAOI21X1_64 OAI21X1_95/Y NAND3X1_93/Y AND2X2_17/Y gnd AOI21X1_64/Y vdd AOI21X1
XAOI21X1_63 OAI21X1_96/Y NAND3X1_95/Y NAND3X1_96/A gnd AOI21X1_63/Y vdd AOI21X1
XNAND3X1_96 NAND3X1_96/A NAND3X1_95/Y OAI21X1_96/Y gnd NAND3X1_96/Y vdd NAND3X1
XNAND2X1_91 A<2> B<4> gnd NAND2X1_91/Y vdd NAND2X1
XNAND2X1_81 A<1> B<4> gnd INVX1_39/A vdd NAND2X1
XNAND3X1_72 B<3> A<2> INVX1_39/A gnd NAND3X1_73/B vdd NAND3X1
XNAND2X1_82 B<3> A<1> gnd OAI21X1_66/C vdd NAND2X1
XOAI21X1_66 gnd INVX2_9/Y OAI21X1_66/C gnd OAI21X1_66/Y vdd OAI21X1
XNOR3X1_7 NOR3X1_7/A NOR3X1_7/B NOR3X1_7/C gnd NOR3X1_7/Y vdd NOR3X1
XOAI21X1_81 NOR3X1_7/B NOR3X1_7/C NOR3X1_7/A gnd OAI21X1_81/Y vdd OAI21X1
XOAI21X1_83 NOR3X1_7/B NOR3X1_7/C vdd gnd OAI21X1_83/Y vdd OAI21X1
XAOI21X1_60 vdd NAND3X1_67/Y vdd gnd AOI21X1_60/Y vdd AOI21X1
XAOI21X1_51 OAI21X1_69/Y NAND3X1_61/Y OAI22X1_5/Y gnd AOI21X1_51/Y vdd AOI21X1
XNAND3X1_62 NAND3X1_61/Y OAI21X1_69/Y OAI22X1_5/Y gnd NAND3X1_62/Y vdd NAND3X1
XINVX1_34 INVX1_34/A gnd INVX1_34/Y vdd INVX1
XNAND2X1_79 INVX1_34/Y XNOR2X1_6/Y gnd NAND2X1_79/Y vdd NAND2X1
XNOR2X1_33 INVX1_34/Y XNOR2X1_6/Y gnd NOR2X1_33/Y vdd NOR2X1
XNAND2X1_80 INVX1_34/A XNOR2X1_7/Y gnd NAND2X1_80/Y vdd NAND2X1
XNOR2X1_32 INVX1_34/A XNOR2X1_7/Y gnd NOR2X1_32/Y vdd NOR2X1
XFILL_8_2 gnd vdd FILL
XFILL_8_1 gnd vdd FILL
XOAI21X1_31 INVX1_9/Y AOI21X1_18/Y NOR2X1_12/B gnd AOI22X1_6/C vdd OAI21X1
XOAI21X1_21 AOI21X1_19/Y AOI21X1_18/Y OAI21X1_7/Y gnd gnd vdd OAI21X1
XOAI21X1_50 AOI21X1_32/Y OAI21X1_41/B OAI22X1_2/C gnd AOI22X1_8/B vdd OAI21X1
XINVX1_15 INVX1_15/A gnd INVX1_15/Y vdd INVX1
XAOI21X1_31 NAND3X1_43/Y OAI21X1_39/Y INVX1_15/Y gnd OAI21X1_41/B vdd AOI21X1
XNAND3X1_46 INVX1_15/Y OAI21X1_39/Y NAND3X1_43/Y gnd NAND3X1_46/Y vdd NAND3X1
XNAND2X1_48 NAND2X1_47/Y AOI21X1_30/Y gnd NAND3X1_45/C vdd NAND2X1
XOAI21X1_43 AOI21X1_30/Y NAND2X1_47/Y OAI21X1_43/C gnd gnd vdd OAI21X1
XNAND3X1_43 OAI21X1_38/Y OR2X2_4/B AOI21X1_30/Y gnd NAND3X1_43/Y vdd NAND3X1
XOAI21X1_7 INVX1_55/Y OAI21X1_7/B INVX1_8/A gnd OAI21X1_7/Y vdd OAI21X1
XNAND3X1_12 INVX1_55/Y OAI21X1_3/Y NAND3X1_9/Y gnd AOI21X1_9/B vdd NAND3X1
XAOI21X1_5 NAND3X1_9/Y OAI21X1_3/Y INVX1_55/Y gnd NOR3X1_3/C vdd AOI21X1
XINVX1_55 INVX1_55/A gnd INVX1_55/Y vdd INVX1
XINVX1_20 INVX1_20/A gnd INVX1_20/Y vdd INVX1
XNAND3X1_42 INVX1_20/Y OAI21X1_44/C NAND3X1_41/Y gnd OR2X2_4/B vdd NAND3X1
XAOI21X1_29 NAND2X1_44/Y vdd INVX1_17/A gnd OAI21X1_38/A vdd AOI21X1
XNAND3X1_40 INVX1_17/A vdd NAND2X1_44/Y gnd OAI21X1_44/C vdd NAND3X1
XOAI21X1_44 INVX1_19/A INVX1_18/A OAI21X1_44/C gnd INVX1_23/A vdd OAI21X1
XBUFX4_4 BUFX4_4/A gnd BUFX4_4/Y vdd BUFX4
XNAND2X1_42 A<5> B<6> gnd INVX1_19/A vdd NAND2X1
XNOR2X1_22 INVX2_2/Y INVX2_3/Y gnd NOR2X1_22/Y vdd NOR2X1
XOAI22X1_4 vdd INVX2_3/Y BUFX4_4/Y INVX2_2/Y gnd OAI22X1_4/Y vdd OAI22X1
XOAI21X1_120 gnd NOR2X1_45/Y OAI21X1_120/C gnd INVX1_55/A vdd OAI21X1
XINVX1_49 gnd gnd INVX1_49/Y vdd INVX1
XNAND3X1_121 INVX1_49/Y OAI21X1_104/Y NAND2X1_110/Y gnd NAND3X1_121/Y vdd NAND3X1
XNAND3X1_106 gnd OAI21X1_104/Y NAND2X1_110/Y gnd NAND3X1_106/Y vdd NAND3X1
XNAND2X1_110 INVX1_50/A NOR2X1_45/B gnd NAND2X1_110/Y vdd NAND2X1
XNOR2X1_45 INVX1_50/A NOR2X1_45/B gnd NOR2X1_45/Y vdd NOR2X1
XNOR2X1_42 vdd BUFX4_4/Y gnd INVX1_50/A vdd NOR2X1
XOAI21X1_104 vdd BUFX4_1/Y NOR2X1_44/B gnd OAI21X1_104/Y vdd OAI21X1
XINVX1_50 INVX1_50/A gnd INVX1_50/Y vdd INVX1
XNOR2X1_44 INVX1_50/Y NOR2X1_44/B gnd NOR2X1_44/Y vdd NOR2X1
XOAI21X1_103 INVX1_43/A NOR2X1_43/Y NAND3X1_87/C gnd NOR2X1_45/B vdd OAI21X1
XAOI22X1_16 NOR2X1_39/Y AND2X2_19/Y INVX1_43/Y OAI21X1_90/Y gnd NOR2X1_44/B vdd AOI22X1
XINVX1_43 INVX1_43/A gnd INVX1_43/Y vdd INVX1
XNAND3X1_87 INVX1_43/Y OAI21X1_90/Y NAND3X1_87/C gnd AND2X2_17/B vdd NAND3X1
XNOR2X1_39 INVX4_1/Y INVX4_4/Y gnd NOR2X1_39/Y vdd NOR2X1
XOAI21X1_90 INVX4_1/Y vdd OAI21X1_90/C gnd OAI21X1_90/Y vdd OAI21X1
XOAI21X1_98 AOI21X1_63/Y AOI21X1_64/Y OAI21X1_89/Y gnd OAI21X1_98/Y vdd OAI21X1
XOAI21X1_97 AOI21X1_63/Y AOI21X1_64/Y AOI21X1_62/Y gnd OAI21X1_97/Y vdd OAI21X1
XOAI21X1_76 INVX4_1/Y INVX4_4/Y INVX1_39/A gnd OAI21X1_77/C vdd OAI21X1
XOAI21X1_77 OAI21X1_66/C NAND2X1_91/Y OAI21X1_77/C gnd OAI21X1_77/Y vdd OAI21X1
XOAI21X1_82 INVX4_1/Y INVX4_4/Y INVX1_39/Y gnd NAND3X1_73/C vdd OAI21X1
XINVX1_39 INVX1_39/A gnd INVX1_39/Y vdd INVX1
XNAND3X1_73 INVX1_41/A NAND3X1_73/B NAND3X1_73/C gnd NAND3X1_73/Y vdd NAND3X1
XNOR2X1_31 INVX4_1/Y gnd gnd INVX2_8/A vdd NOR2X1
XOAI21X1_67 INVX1_39/A INVX2_8/Y OAI21X1_66/Y gnd OR2X2_7/B vdd OAI21X1
XAOI21X1_62 AOI21X1_62/A OAI21X1_81/Y NOR3X1_7/Y gnd AOI21X1_62/Y vdd AOI21X1
XOAI21X1_89 AOI21X1_60/Y OAI21X1_89/B OAI21X1_89/C gnd OAI21X1_89/Y vdd OAI21X1
XNAND3X1_74 NAND3X1_67/Y vdd NOR3X1_7/A gnd NAND3X1_74/Y vdd NAND3X1
XNAND3X1_69 NAND3X1_67/Y vdd vdd gnd NAND3X1_69/Y vdd NAND3X1
XOAI21X1_75 OR2X2_7/B AOI21X1_51/Y NAND3X1_62/Y gnd OAI21X1_75/Y vdd OAI21X1
XINVX2_8 INVX2_8/A gnd INVX2_8/Y vdd INVX2
XNAND3X1_58 INVX2_8/Y NAND2X1_80/Y NAND2X1_79/Y gnd NAND3X1_58/Y vdd NAND3X1
XOAI21X1_63 NOR2X1_32/Y NOR2X1_33/Y INVX2_8/A gnd OAI21X1_63/Y vdd OAI21X1
XNAND3X1_59 INVX2_8/A NAND2X1_80/Y NAND2X1_79/Y gnd NAND3X1_59/Y vdd NAND3X1
XOAI21X1_65 INVX2_8/Y NOR2X1_33/Y NAND2X1_79/Y gnd OAI21X1_65/Y vdd OAI21X1
XOAI21X1_64 NOR2X1_32/Y NOR2X1_33/Y INVX2_8/Y gnd OAI21X1_64/Y vdd OAI21X1
XAOI22X1_6 AOI22X1_6/A AOI22X1_6/B AOI22X1_6/C AOI22X1_6/D gnd AOI22X1_6/Y vdd AOI22X1
XOAI22X1_2 NOR2X1_12/A NOR2X1_12/B OAI22X1_2/C OAI22X1_2/D gnd OAI22X1_2/Y vdd OAI22X1
XNAND3X1_47 OAI21X1_43/C NAND3X1_46/Y OAI22X1_2/C gnd AOI22X1_6/B vdd NAND3X1
XNAND2X1_57 OAI21X1_43/C NAND3X1_46/Y gnd OAI22X1_2/D vdd NAND2X1
XNAND2X1_61 NAND3X1_25/Y NAND3X1_27/Y gnd NOR2X1_19/B vdd NAND2X1
XAOI21X1_36 NAND3X1_25/Y NAND3X1_27/Y AOI21X1_20/Y gnd OAI22X1_3/A vdd AOI21X1
XNAND3X1_29 NAND3X1_25/Y NAND3X1_27/Y AOI21X1_20/Y gnd AOI22X1_4/A vdd NAND3X1
XAOI22X1_4 AOI22X1_4/A gnd AOI22X1_4/C AOI22X1_4/D gnd AND2X2_6/A vdd AOI22X1
XINVX1_8 INVX1_8/A gnd INVX1_8/Y vdd INVX1
XAOI21X1_20 INVX1_55/A OAI21X1_4/Y INVX1_8/Y gnd AOI21X1_20/Y vdd AOI21X1
XNAND3X1_13 AOI21X1_9/A AOI21X1_9/B AOI21X1_7/Y gnd AOI22X1_4/D vdd NAND3X1
XNAND3X1_11 INVX1_55/A INVX1_8/A OAI21X1_4/Y gnd AOI21X1_9/A vdd NAND3X1
XNAND2X1_10 AOI22X1_4/C AOI22X1_4/D gnd XOR2X1_1/B vdd NAND2X1
XAOI21X1_6 OAI21X1_4/Y INVX1_8/A INVX1_55/A gnd NOR3X1_3/B vdd AOI21X1
XBUFX4_3 BUFX4_4/A gnd BUFX4_3/Y vdd BUFX4
XBUFX4_2 BUFX4_4/A gnd BUFX4_2/Y vdd BUFX4
XINVX8_1 B<6> gnd BUFX4_4/A vdd INVX8
XBUFX4_1 BUFX4_4/A gnd BUFX4_1/Y vdd BUFX4
XNOR2X1_21 vdd BUFX4_3/Y gnd NOR2X1_21/Y vdd NOR2X1
XOAI21X1_57 vdd BUFX4_1/Y NOR2X1_22/Y gnd XOR2X1_4/B vdd OAI21X1
XNAND2X1_53 OR2X2_6/A OAI21X1_48/Y gnd OR2X2_4/A vdd NAND2X1
XNAND2X1_63 OAI22X1_4/Y NAND2X1_63/B gnd OR2X2_6/B vdd NAND2X1
XOAI21X1_113 NOR2X1_44/Y NOR2X1_45/Y gnd gnd NAND2X1_120/B vdd OAI21X1
XNAND2X1_120 NAND3X1_121/Y NAND2X1_120/B gnd AOI21X1_74/C vdd NAND2X1
XOAI21X1_105 NOR2X1_44/Y NOR2X1_45/Y INVX1_49/Y gnd NAND2X1_111/B vdd OAI21X1
XNAND2X1_111 NAND3X1_106/Y NAND2X1_111/B gnd AOI21X1_4/A vdd NAND2X1
XAOI21X1_75 AOI21X1_4/B AOI21X1_75/B AOI21X1_4/A gnd AOI21X1_75/Y vdd AOI21X1
XNAND3X1_120 AOI21X1_4/A AOI21X1_75/B AOI21X1_4/B gnd AOI21X1_80/B vdd NAND3X1
XNAND3X1_123 AOI21X1_74/C AOI21X1_74/B AOI21X1_74/A gnd AOI21X1_80/A vdd NAND3X1
XAOI21X1_74 AOI21X1_74/A AOI21X1_74/B AOI21X1_74/C gnd vdd vdd AOI21X1
XNOR2X1_41 gnd BUFX4_3/Y gnd NOR2X1_41/Y vdd NOR2X1
XOAI21X1_88 gnd BUFX4_2/Y OAI21X1_88/C gnd OAI21X1_88/Y vdd OAI21X1
XNAND2X1_108 NOR2X1_41/Y OAI21X1_87/Y gnd INVX1_48/A vdd NAND2X1
XOAI21X1_102 INVX1_46/Y AOI21X1_68/Y INVX1_54/A gnd AOI21X1_80/C vdd OAI21X1
XAOI21X1_68 NAND3X1_94/Y NAND3X1_96/Y OAI21X1_89/Y gnd AOI21X1_68/Y vdd AOI21X1
XNAND3X1_97 NAND3X1_94/Y NAND3X1_96/Y OAI21X1_89/Y gnd INVX1_54/A vdd NAND3X1
XNAND3X1_99 NAND3X1_94/Y NAND3X1_96/Y AOI21X1_62/Y gnd NAND3X1_99/Y vdd NAND3X1
XOAI21X1_87 INVX1_41/A OAI21X1_77/Y NAND3X1_66/C gnd OAI21X1_87/Y vdd OAI21X1
XNAND2X1_90 INVX1_39/Y NOR2X1_39/Y gnd NAND3X1_66/C vdd NAND2X1
XNAND3X1_66 INVX1_41/A OAI21X1_77/C NAND3X1_66/C gnd AOI22X1_11/A vdd NAND3X1
XNAND2X1_92 INVX1_41/Y OAI21X1_77/Y gnd AOI22X1_11/B vdd NAND2X1
XNAND2X1_88 INVX1_39/Y INVX2_8/A gnd INVX1_40/A vdd NAND2X1
XNAND2X1_93 AOI22X1_11/A AOI22X1_11/B gnd AOI21X1_62/A vdd NAND2X1
XAOI22X1_11 AOI22X1_11/A AOI22X1_11/B NAND3X1_74/Y OAI21X1_83/Y gnd NOR3X1_8/A vdd
+ AOI22X1
XNAND3X1_75 NAND3X1_74/Y OAI21X1_89/B OAI21X1_83/Y gnd NAND3X1_75/Y vdd NAND3X1
XNAND3X1_70 NAND3X1_69/Y OAI21X1_81/Y AOI21X1_62/A gnd NAND3X1_78/A vdd NAND3X1
XAOI21X1_55 OAI21X1_81/Y NAND3X1_69/Y AOI21X1_62/A gnd NOR3X1_8/B vdd AOI21X1
XINVX1_37 OR2X2_7/B gnd INVX1_37/Y vdd INVX1
XNAND2X1_87 NAND3X1_62/Y OAI21X1_72/Y gnd OR2X2_7/A vdd NAND2X1
XAOI21X1_47 OAI21X1_72/Y NAND3X1_62/Y INVX1_37/Y gnd INVX1_38/A vdd AOI21X1
XAOI21X1_54 INVX1_37/Y OAI21X1_72/Y NOR3X1_5/Y gnd vdd vdd AOI21X1
XINVX1_33 INVX1_33/A gnd INVX1_33/Y vdd INVX1
XAOI21X1_42 OAI21X1_63/Y NAND3X1_58/Y INVX1_33/Y gnd NOR2X1_34/A vdd AOI21X1
XAOI21X1_48 NAND2X1_80/Y INVX2_8/A NOR2X1_32/Y gnd NOR3X1_6/C vdd AOI21X1
XAOI21X1_43 OAI21X1_64/Y NAND3X1_59/Y INVX1_33/A gnd NOR2X1_34/B vdd AOI21X1
XNAND3X1_60 INVX1_33/A NAND3X1_59/Y OAI21X1_64/Y gnd NAND3X1_60/Y vdd NAND3X1
XBUFX2_4 BUFX2_4/A gnd S<3> vdd BUFX2
XFILL_10_1 gnd vdd FILL
XINVX1_13 INVX1_13/A gnd INVX1_13/Y vdd INVX1
XNAND3X1_48 AOI22X1_6/A AOI22X1_6/B NAND3X1_48/C gnd NAND3X1_48/Y vdd NAND3X1
XNAND2X1_49 AOI22X1_6/B AOI22X1_6/A gnd NAND3X1_49/B vdd NAND2X1
XNAND2X1_58 AOI22X1_8/B OAI22X1_2/Y gnd NAND2X1_58/Y vdd NAND2X1
XNAND3X1_28 NAND3X1_25/Y NAND3X1_27/Y OAI21X1_7/Y gnd NAND3X1_28/Y vdd NAND3X1
XAOI21X1_17 NAND3X1_27/Y NAND3X1_25/Y OAI21X1_7/Y gnd INVX1_7/A vdd AOI21X1
XAOI22X1_8 OAI22X1_2/Y AOI22X1_8/B INVX1_7/Y AOI22X1_8/D gnd AOI22X1_8/Y vdd AOI22X1
XOAI21X1_51 AOI21X1_20/Y NOR2X1_19/B OAI21X1_6/C gnd AOI22X1_8/D vdd OAI21X1
XNOR2X1_19 OAI21X1_7/Y NOR2X1_19/B gnd OAI22X1_3/B vdd NOR2X1
XOAI22X1_3 OAI22X1_3/A OAI22X1_3/B NOR2X1_2/A NOR3X1_3/Y gnd OAI22X1_3/Y vdd OAI22X1
XNOR2X1_2 NOR2X1_2/A NOR3X1_3/Y gnd NOR2X1_2/Y vdd NOR2X1
XAOI21X1_9 AOI21X1_9/A AOI21X1_9/B AOI21X1_7/Y gnd NOR2X1_2/A vdd AOI21X1
XNAND3X1_14 AOI21X1_9/A AOI21X1_9/B NOR3X1_3/A gnd OAI21X1_6/C vdd NAND3X1
XOAI21X1_5 NOR3X1_3/B NOR3X1_3/C NOR3X1_3/A gnd AOI22X1_4/C vdd OAI21X1
XNOR3X1_3 NOR3X1_3/A NOR3X1_3/B NOR3X1_3/C gnd NOR3X1_3/Y vdd NOR3X1
XXOR2X1_1 XOR2X1_1/A XOR2X1_1/B gnd XOR2X1_1/Y vdd XOR2X1
XOR2X2_4 OR2X2_4/A OR2X2_4/B gnd OR2X2_4/Y vdd OR2X2
XDFFPOSX1_12 BUFX2_9/A clk XOR2X1_1/Y gnd vdd DFFPOSX1
XNAND2X1_62 NOR2X1_21/Y NOR2X1_22/Y gnd NAND2X1_63/B vdd NAND2X1
XNAND2X1_64 OR2X2_6/B OR2X2_6/A gnd NAND2X1_64/Y vdd NAND2X1
XOR2X2_6 OR2X2_6/A OR2X2_6/B gnd OR2X2_6/Y vdd OR2X2
XAOI21X1_7 INVX1_48/Y AOI21X1_7/B INVX1_1/Y gnd AOI21X1_7/Y vdd AOI21X1
XINVX1_1 INVX1_1/A gnd INVX1_1/Y vdd INVX1
XOAI21X1_119 INVX1_48/A AOI21X1_80/Y INVX1_1/A gnd NOR3X1_3/A vdd OAI21X1
XAOI21X1_80 AOI21X1_80/A AOI21X1_80/B AOI21X1_80/C gnd AOI21X1_80/Y vdd AOI21X1
XNAND3X1_124 AOI21X1_80/B AOI21X1_80/C AOI21X1_80/A gnd INVX1_1/A vdd NAND3X1
XNAND3X1_126 AOI21X1_80/B AOI21X1_80/A AOI21X1_73/Y gnd AOI21X1_76/A vdd NAND3X1
XINVX2_6 A<0> gnd gnd vdd INVX2
XINVX1_54 INVX1_54/A gnd INVX1_54/Y vdd INVX1
XAOI21X1_73 INVX1_46/A OAI21X1_97/Y INVX1_54/Y gnd AOI21X1_73/Y vdd AOI21X1
XINVX1_46 INVX1_46/A gnd INVX1_46/Y vdd INVX1
XNAND2X1_99 NAND3X1_86/Y OAI21X1_88/Y gnd INVX1_46/A vdd NAND2X1
XAOI22X1_15 OAI21X1_88/Y NAND3X1_86/Y NAND3X1_99/Y OAI21X1_98/Y gnd NOR2X1_46/A vdd
+ AOI22X1
XNAND3X1_100 INVX1_46/Y NAND3X1_99/Y OAI21X1_98/Y gnd NAND3X1_100/Y vdd NAND3X1
XAOI21X1_66 OAI21X1_97/Y INVX1_54/A INVX1_46/A gnd NOR2X1_46/B vdd AOI21X1
XNAND3X1_98 INVX1_46/A INVX1_54/A OAI21X1_97/Y gnd NAND3X1_98/Y vdd NAND3X1
XNAND3X1_86 NAND3X1_66/C NOR2X1_41/Y NAND2X1_98/B gnd NAND3X1_86/Y vdd NAND3X1
XNAND3X1_71 INVX1_41/Y OAI21X1_77/C NAND3X1_66/C gnd NAND2X1_98/B vdd NAND3X1
XINVX1_41 INVX1_41/A gnd INVX1_41/Y vdd INVX1
XNAND2X1_98 NAND3X1_73/Y NAND2X1_98/B gnd OAI21X1_89/B vdd NAND2X1
XOAI21X1_86 INVX1_40/A AOI21X1_59/Y NAND3X1_76/Y gnd OAI21X1_86/Y vdd OAI21X1
XAOI21X1_59 NAND3X1_78/A NAND3X1_75/Y OAI21X1_75/Y gnd AOI21X1_59/Y vdd AOI21X1
XNAND3X1_76 NAND3X1_75/Y NAND3X1_78/A OAI21X1_75/Y gnd NAND3X1_76/Y vdd NAND3X1
XNAND3X1_78 NAND3X1_78/A NAND3X1_75/Y vdd gnd NAND3X1_78/Y vdd NAND3X1
XOAI21X1_85 NOR3X1_8/A NOR3X1_8/B OAI21X1_75/Y gnd OAI21X1_85/Y vdd OAI21X1
XNOR2X1_37 OR2X2_7/B OR2X2_7/A gnd NOR3X1_6/A vdd NOR2X1
XOR2X2_7 OR2X2_7/A OR2X2_7/B gnd OR2X2_7/Y vdd OR2X2
XINVX1_38 INVX1_38/A gnd INVX1_38/Y vdd INVX1
XNAND3X1_64 OR2X2_7/Y INVX1_38/Y OAI21X1_65/Y gnd NAND3X1_64/Y vdd NAND3X1
XNAND3X1_63 INVX1_38/Y OR2X2_7/Y NOR3X1_6/C gnd NAND3X1_63/Y vdd NAND3X1
XNOR2X1_34 NOR2X1_34/A NOR2X1_34/B gnd NOR2X1_34/Y vdd NOR2X1
XDFFPOSX1_7 BUFX2_4/A clk NOR2X1_34/Y gnd vdd DFFPOSX1
XFILL_11_1 gnd vdd FILL
XINVX1_14 INVX1_14/A gnd INVX1_14/Y vdd INVX1
XOAI21X1_32 INVX1_14/Y XNOR2X1_2/A INVX1_13/Y gnd NAND3X1_48/C vdd OAI21X1
XNAND2X1_59 NAND3X1_49/B INVX1_14/A gnd NAND2X1_60/B vdd NAND2X1
XNAND2X1_60 NAND2X1_58/Y NAND2X1_60/B gnd NAND2X1_60/Y vdd NAND2X1
XAOI22X1_7 AOI22X1_8/B OAI22X1_2/Y AOI22X1_7/C AOI22X1_6/Y gnd AOI22X1_7/Y vdd AOI22X1
XOAI21X1_22 INVX1_7/A OAI21X1_6/C NAND3X1_28/Y gnd AOI22X1_7/C vdd OAI21X1
XINVX1_7 INVX1_7/A gnd INVX1_7/Y vdd INVX1
XNAND2X1_27 NAND3X1_28/Y INVX1_7/Y gnd XNOR2X1_1/B vdd NAND2X1
XNAND3X1_52 AOI22X1_6/Y XOR2X1_1/A AND2X2_6/A gnd AOI21X1_40/A vdd NAND3X1
XOAI21X1_52 OAI21X1_6/B OAI22X1_3/Y AOI22X1_8/Y gnd OAI21X1_52/Y vdd OAI21X1
XOAI21X1_6 NOR2X1_2/Y OAI21X1_6/B OAI21X1_6/C gnd OAI21X1_6/Y vdd OAI21X1
XAOI21X1_35 AOI21X1_40/A AOI22X1_7/Y NAND2X1_56/Y gnd NOR2X1_20/A vdd AOI21X1
XAOI21X1_40 AOI21X1_40/A AOI22X1_7/Y NAND3X1_57/Y gnd AOI21X1_40/Y vdd AOI21X1
XNAND2X1_56 INVX1_24/Y OR2X2_5/Y gnd NAND2X1_56/Y vdd NAND2X1
XNAND3X1_57 INVX1_24/Y AND2X2_8/Y OR2X2_5/Y gnd NAND3X1_57/Y vdd NAND3X1
XINVX1_24 INVX1_24/A gnd INVX1_24/Y vdd INVX1
XAOI21X1_34 OAI21X1_49/Y NAND3X1_51/Y gnd gnd INVX1_24/A vdd AOI21X1
XNAND2X1_55 NAND3X1_51/Y OAI21X1_49/Y gnd OR2X2_5/A vdd NAND2X1
XNAND3X1_51 INVX1_23/A AOI21X1_38/B OR2X2_4/Y gnd NAND3X1_51/Y vdd NAND3X1
XAND2X2_7 OR2X2_4/A OR2X2_4/B gnd AND2X2_7/Y vdd AND2X2
XOAI21X1_53 INVX1_23/Y AND2X2_7/Y OR2X2_4/Y gnd NAND2X1_66/A vdd OAI21X1
XOAI21X1_49 NOR2X1_16/Y AND2X2_7/Y INVX1_23/Y gnd OAI21X1_49/Y vdd OAI21X1
XINVX1_23 INVX1_23/A gnd INVX1_23/Y vdd INVX1
XNAND2X1_54 OR2X2_4/B OR2X2_4/A gnd AOI21X1_38/B vdd NAND2X1
XNOR2X1_16 OR2X2_4/B OR2X2_4/A gnd NOR2X1_16/Y vdd NOR2X1
XAOI21X1_38 INVX1_23/A AOI21X1_38/B NOR2X1_16/Y gnd AOI21X1_38/Y vdd AOI21X1
XNAND2X1_66 NAND2X1_66/A XNOR2X1_3/Y gnd AND2X2_8/B vdd NAND2X1
XAOI21X1_41 NOR2X1_21/Y NOR2X1_22/Y NOR2X1_23/Y gnd AOI21X1_41/Y vdd AOI21X1
XXOR2X1_3 XOR2X1_3/A XOR2X1_3/B gnd XOR2X1_3/Y vdd XOR2X1
XNAND2X1_65 NAND2X1_64/Y OR2X2_6/Y gnd XOR2X1_3/A vdd NAND2X1
XXNOR2X1_3 XNOR2X1_3/A XOR2X1_3/B gnd XNOR2X1_3/Y vdd XNOR2X1
XNAND3X1_125 INVX1_48/Y INVX1_1/A AOI21X1_7/B gnd AOI22X1_21/C vdd NAND3X1
XINVX1_48 INVX1_48/A gnd INVX1_48/Y vdd INVX1
XOAI21X1_115 vdd AOI21X1_75/Y AOI21X1_73/Y gnd AOI21X1_7/B vdd OAI21X1
XOAI21X1_116 vdd AOI21X1_75/Y AOI21X1_80/C gnd AOI21X1_76/B vdd OAI21X1
XAOI21X1_76 AOI21X1_76/A AOI21X1_76/B INVX1_48/A gnd AOI21X1_76/Y vdd AOI21X1
XNAND3X1_127 INVX1_48/A AOI21X1_76/B AOI21X1_76/A gnd AOI22X1_21/D vdd NAND3X1
XINVX1_47 INVX1_47/A gnd INVX1_47/Y vdd INVX1
XNAND3X1_128 INVX1_47/Y AOI22X1_21/C AOI22X1_21/D gnd INVX1_2/A vdd NAND3X1
XAOI22X1_21 OAI21X1_86/Y NOR2X1_46/Y AOI22X1_21/C AOI22X1_21/D gnd AOI22X1_21/Y vdd
+ AOI22X1
XNOR2X1_46 NOR2X1_46/A NOR2X1_46/B gnd NOR2X1_46/Y vdd NOR2X1
XNAND3X1_101 NAND3X1_98/Y NAND3X1_100/Y OAI21X1_86/Y gnd INVX1_47/A vdd NAND3X1
XNAND3X1_103 NAND3X1_98/Y NAND3X1_100/Y AOI21X1_65/Y gnd AOI21X1_78/A vdd NAND3X1
XOAI21X1_99 NOR2X1_46/A NOR2X1_46/B AOI21X1_65/Y gnd OAI21X1_99/Y vdd OAI21X1
XOAI21X1_100 NOR2X1_46/A NOR2X1_46/B OAI21X1_100/C gnd AOI21X1_78/B vdd OAI21X1
XNAND3X1_104 AOI21X1_78/C AOI21X1_78/B AOI21X1_78/A gnd AOI21X1_79/A vdd NAND3X1
XAOI21X1_78 AOI21X1_78/A AOI21X1_78/B AOI21X1_78/C gnd AOI21X1_78/Y vdd AOI21X1
XAOI21X1_65 INVX1_40/Y OAI21X1_84/Y NOR3X1_8/Y gnd AOI21X1_65/Y vdd AOI21X1
XOAI21X1_84 NOR3X1_8/A NOR3X1_8/B vdd gnd OAI21X1_84/Y vdd OAI21X1
XNOR3X1_8 NOR3X1_8/A NOR3X1_8/B vdd gnd NOR3X1_8/Y vdd NOR3X1
XOAI21X1_74 NOR3X1_6/A INVX1_38/A NOR3X1_6/C gnd OAI21X1_74/Y vdd OAI21X1
XNOR3X1_6 NOR3X1_6/A INVX1_38/A NOR3X1_6/C gnd NOR3X1_6/Y vdd NOR3X1
XOAI21X1_73 NOR3X1_6/A INVX1_38/A OAI21X1_65/Y gnd AOI21X1_49/A vdd OAI21X1
XAOI21X1_49 AOI21X1_49/A NAND3X1_63/Y NAND3X1_60/Y gnd NOR2X1_38/A vdd AOI21X1
XFILL_12_3 gnd vdd FILL
XFILL_12_2 gnd vdd FILL
XFILL_12_1 gnd vdd FILL
XDFFPOSX1_14 BUFX2_11/A clk XNOR2X1_2/Y gnd vdd DFFPOSX1
XOAI21X1_42 AOI22X1_7/C AND2X2_6/Y INVX1_14/A gnd NAND3X1_49/C vdd OAI21X1
XAOI21X1_21 AND2X2_6/A XOR2X1_1/A AOI22X1_7/C gnd XNOR2X1_2/A vdd AOI21X1
XAND2X2_6 AND2X2_6/A XOR2X1_1/A gnd AND2X2_6/Y vdd AND2X2
XXNOR2X1_1 OAI21X1_6/Y XNOR2X1_1/B gnd XNOR2X1_1/Y vdd XNOR2X1
XAOI21X1_37 OAI21X1_52/Y NAND2X1_60/Y NOR2X1_18/Y gnd NOR2X1_20/B vdd AOI21X1
XNOR2X1_20 NOR2X1_20/A NOR2X1_20/B gnd NOR2X1_20/Y vdd NOR2X1
XNAND3X1_53 NOR2X1_18/Y NAND2X1_60/Y OAI21X1_52/Y gnd NAND3X1_54/C vdd NAND3X1
XNAND3X1_55 NAND2X1_60/Y NOR3X1_4/Y OAI21X1_52/Y gnd NAND3X1_55/Y vdd NAND3X1
XNAND3X1_54 OR2X2_5/Y AND2X2_8/Y NAND3X1_54/C gnd NAND3X1_54/Y vdd NAND3X1
XNOR2X1_18 INVX1_24/A NOR3X1_4/C gnd NOR2X1_18/Y vdd NOR2X1
XOAI21X1_55 NOR3X1_4/C NOR2X1_20/A NOR3X1_4/B gnd OAI21X1_55/Y vdd OAI21X1
XNOR3X1_4 INVX1_24/A NOR3X1_4/B NOR3X1_4/C gnd NOR3X1_4/Y vdd NOR3X1
XNOR2X1_17 OR2X2_5/B OR2X2_5/A gnd NOR3X1_4/C vdd NOR2X1
XINVX1_25 gnd gnd OR2X2_5/B vdd INVX1
XOR2X2_5 OR2X2_5/A OR2X2_5/B gnd OR2X2_5/Y vdd OR2X2
XOAI21X1_56 NOR3X1_4/B OR2X2_5/Y AND2X2_8/B gnd INVX1_26/A vdd OAI21X1
XAND2X2_8 AND2X2_8/A AND2X2_8/B gnd AND2X2_8/Y vdd AND2X2
XNAND2X1_68 AND2X2_8/B AND2X2_8/A gnd NOR3X1_4/B vdd NAND2X1
XNAND2X1_67 AOI21X1_38/Y XOR2X1_3/Y gnd AND2X2_8/A vdd NAND2X1
XXOR2X1_4 XOR2X1_4/A XOR2X1_4/B gnd XOR2X1_4/Y vdd XOR2X1
XNOR2X1_23 XOR2X1_4/B XOR2X1_4/A gnd NOR2X1_23/Y vdd NOR2X1
XINVX1_27 OR2X2_6/Y gnd INVX1_27/Y vdd INVX1
XAOI21X1_39 XOR2X1_3/B NAND2X1_64/Y INVX1_27/Y gnd XOR2X1_4/A vdd AOI21X1
XAOI21X1_77 AOI21X1_7/B INVX1_1/A INVX1_48/Y gnd AOI21X1_77/Y vdd AOI21X1
XAOI21X1_8 AOI21X1_8/A AOI21X1_8/B INVX1_2/Y gnd OAI21X1_6/B vdd AOI21X1
XINVX1_2 INVX1_2/A gnd INVX1_2/Y vdd INVX1
XOAI21X1_117 AOI21X1_77/Y AOI21X1_76/Y INVX1_47/A gnd AOI21X1_8/B vdd OAI21X1
XNAND2X1_121 INVX1_2/A AOI21X1_8/B gnd XNOR2X1_9/A vdd NAND2X1
XOAI21X1_118 AOI22X1_21/Y AOI21X1_79/Y INVX1_2/A gnd XOR2X1_1/A vdd OAI21X1
XAOI21X1_67 OAI21X1_99/Y INVX1_47/A AOI21X1_58/Y gnd AOI21X1_67/Y vdd AOI21X1
XOAI21X1_101 OAI21X1_101/A AOI21X1_67/Y OAI21X1_101/C gnd AOI21X1_8/A vdd OAI21X1
XNAND3X1_102 INVX1_47/A AOI21X1_58/Y OAI21X1_99/Y gnd NAND2X1_107/A vdd NAND3X1
XNAND2X1_107 NAND2X1_107/A AOI21X1_79/A gnd XNOR2X1_8/A vdd NAND2X1
XXNOR2X1_8 XNOR2X1_8/A XNOR2X1_8/B gnd XNOR2X1_8/Y vdd XNOR2X1
XAOI21X1_79 AOI21X1_79/A XNOR2X1_8/B AOI21X1_78/Y gnd AOI21X1_79/Y vdd AOI21X1
XNAND3X1_77 INVX1_40/Y NAND3X1_76/Y OAI21X1_84/Y gnd NAND3X1_77/Y vdd NAND3X1
XINVX1_40 INVX1_40/A gnd INVX1_40/Y vdd INVX1
XNAND3X1_81 INVX1_40/A NAND3X1_76/Y OAI21X1_84/Y gnd NAND3X1_83/A vdd NAND3X1
XNAND3X1_79 INVX1_40/A NAND3X1_78/Y OAI21X1_85/Y gnd NAND3X1_79/Y vdd NAND3X1
XNAND3X1_82 INVX1_40/Y NAND3X1_78/Y OAI21X1_85/Y gnd NAND3X1_83/B vdd NAND3X1
XAOI21X1_58 NAND3X1_83/B NAND3X1_83/A NAND3X1_64/Y gnd AOI21X1_58/Y vdd AOI21X1
XNAND3X1_85 NAND3X1_83/A NAND3X1_64/Y NAND3X1_83/B gnd vdd vdd NAND3X1
XNAND3X1_83 NAND3X1_83/A NAND3X1_83/B NOR3X1_6/Y gnd AOI21X1_56/A vdd NAND3X1
XAOI21X1_56 AOI21X1_56/A AOI21X1_56/B NAND3X1_65/Y gnd XNOR2X1_8/B vdd AOI21X1
XAOI21X1_50 NAND3X1_64/Y OAI21X1_74/Y NOR2X1_34/A gnd NOR2X1_38/B vdd AOI21X1
XNAND3X1_65 OAI21X1_74/Y NAND3X1_64/Y NOR2X1_34/A gnd NAND3X1_65/Y vdd NAND3X1
XDFFPOSX1_10 BUFX2_7/A clk XNOR2X1_8/Y gnd vdd DFFPOSX1
XBUFX2_7 BUFX2_7/A gnd S<6> vdd BUFX2
XFILL_13_3 gnd vdd FILL
XFILL_13_2 gnd vdd FILL
XFILL_13_1 gnd vdd FILL
XXNOR2X1_2 XNOR2X1_2/A INVX1_14/A gnd XNOR2X1_2/Y vdd XNOR2X1
XINVX1_6 INVX1_6/A gnd INVX1_6/Y vdd INVX1
XNAND3X1_26 NAND3X1_24/A NAND3X1_24/B AOI21X1_14/Y gnd NAND3X1_27/C vdd NAND3X1
XNAND2X1_50 NAND3X1_49/Y NAND3X1_48/Y gnd NAND2X1_50/Y vdd NAND2X1
XBUFX2_12 BUFX2_12/A gnd S<11> vdd BUFX2
XDFFPOSX1_15 BUFX2_12/A clk NAND2X1_50/Y gnd vdd DFFPOSX1
XBUFX2_13 BUFX2_13/A gnd S<12> vdd BUFX2
XDFFPOSX1_16 BUFX2_13/A clk NOR2X1_20/Y gnd vdd DFFPOSX1
XBUFX2_14 BUFX2_14/A gnd S<13> vdd BUFX2
XNAND2X1_69 OAI21X1_55/Y NAND3X1_54/Y gnd DFFPOSX1_1/D vdd NAND2X1
XDFFPOSX1_1 BUFX2_14/A clk DFFPOSX1_1/D gnd vdd DFFPOSX1
XBUFX2_15 BUFX2_15/A gnd S<14> vdd BUFX2
XDFFPOSX1_2 BUFX2_15/A clk NAND2X1_70/Y gnd vdd DFFPOSX1
XNAND3X1_56 INVX1_26/Y XOR2X1_4/Y NAND3X1_55/Y gnd NAND2X1_70/B vdd NAND3X1
XINVX1_26 INVX1_26/A gnd INVX1_26/Y vdd INVX1
XNAND2X1_70 OAI21X1_58/Y NAND2X1_70/B gnd NAND2X1_70/Y vdd NAND2X1
XOAI21X1_58 INVX1_26/A AOI21X1_40/Y OAI21X1_58/C gnd OAI21X1_58/Y vdd OAI21X1
XINVX1_28 XOR2X1_4/Y gnd INVX1_28/Y vdd INVX1
XOAI21X1_59 INVX1_26/A AOI21X1_40/Y XOR2X1_4/Y gnd vdd vdd OAI21X1
XBUFX2_9 BUFX2_9/A gnd S<8> vdd BUFX2
XDFFPOSX1_13 BUFX2_10/A clk XNOR2X1_1/Y gnd vdd DFFPOSX1
XBUFX2_10 BUFX2_10/A gnd S<9> vdd BUFX2
XNAND2X1_71 AOI21X1_41/Y vdd gnd DFFPOSX1_3/D vdd NAND2X1
XDFFPOSX1_3 BUFX2_16/A DFFPOSX1_3/CLK DFFPOSX1_3/D gnd vdd DFFPOSX1
XBUFX2_16 BUFX2_16/A gnd S<15> vdd BUFX2
XXNOR2X1_9 XNOR2X1_9/A AOI21X1_8/A gnd XNOR2X1_9/Y vdd XNOR2X1
XBUFX2_8 BUFX2_8/A gnd S<7> vdd BUFX2
XDFFPOSX1_11 BUFX2_8/A clk XNOR2X1_9/Y gnd vdd DFFPOSX1
XBUFX2_5 BUFX2_5/A gnd S<4> vdd BUFX2
XDFFPOSX1_8 BUFX2_5/A clk NOR2X1_38/Y gnd vdd DFFPOSX1
XNAND3X1_105 NOR2X1_38/A vdd AOI21X1_78/C gnd OAI21X1_101/A vdd NAND3X1
XNOR2X1_38 NOR2X1_38/A NOR2X1_38/B gnd NOR2X1_38/Y vdd NOR2X1
XNAND3X1_84 NAND3X1_77/Y NAND3X1_79/Y NOR3X1_6/Y gnd AOI21X1_78/C vdd NAND3X1
XNAND3X1_80 NAND3X1_77/Y NAND3X1_64/Y NAND3X1_79/Y gnd AOI21X1_56/B vdd NAND3X1
XAOI21X1_57 AOI21X1_78/C vdd NOR2X1_38/A gnd NOR2X1_40/B vdd AOI21X1
XNOR2X1_40 XNOR2X1_8/B NOR2X1_40/B gnd NOR2X1_40/Y vdd NOR2X1
XDFFPOSX1_9 BUFX2_6/A clk NOR2X1_40/Y gnd vdd DFFPOSX1
XBUFX2_6 BUFX2_6/A gnd S<5> vdd BUFX2
C123 NAND3X1_64/Y 0 2.36fF
C124 NAND3X1_77/Y 0 2.00fF
C125 AOI21X1_78/C 0 3.04fF
C126 XNOR2X1_9/A 0 2.30fF
C127 XNOR2X1_9/Y 0 2.19fF
C128 XNOR2X1_1/Y 0 2.21fF
C129 clk 0 14.18fF
C130 NAND3X1_49/Y 0 2.74fF
C131 XNOR2X1_2/A 0 2.55fF
C132 XNOR2X1_2/Y 0 2.18fF
C133 NAND3X1_83/B 0 2.44fF
C134 NAND3X1_78/Y 0 2.05fF
C135 NAND3X1_76/Y 0 2.16fF
C136 AOI21X1_58/Y 0 2.22fF
C137 OAI21X1_99/Y 0 2.18fF
C138 INVX1_47/A 0 3.08fF
C139 INVX1_2/A 0 2.20fF
C140 INVX1_48/Y 0 2.44fF
C141 INVX1_1/A 0 2.06fF
C142 AOI21X1_7/B 0 2.54fF
C143 NOR3X1_4/B 0 2.46fF
C144 AND2X2_8/Y 0 2.07fF
C145 OR2X2_5/Y 0 2.65fF
C146 OAI21X1_52/Y 0 2.04fF
C147 AND2X2_6/A 0 2.24fF
C148 AOI22X1_7/C 0 2.05fF
C149 vdd 0 565.97fF
C150 NAND3X1_60/Y 0 2.05fF
C151 NOR3X1_8/A 0 2.08fF
C152 NOR3X1_8/B 0 2.14fF
C153 AOI21X1_65/Y 0 2.02fF
C154 NAND3X1_98/Y 0 2.01fF
C155 AOI22X1_21/D 0 2.28fF
C156 AOI21X1_76/A 0 2.02fF
C157 XNOR2X1_3/Y 0 2.09fF
C158 OR2X2_4/A 0 2.04fF
C159 NAND3X1_51/Y 0 2.09fF
C160 OAI21X1_49/Y 0 2.06fF
C161 NAND3X1_75/Y 0 2.41fF
C162 NAND3X1_66/C 0 2.24fF
C163 NAND3X1_86/Y 0 2.02fF
C164 INVX1_54/A 0 2.42fF
C165 AOI21X1_7/Y 0 2.17fF
C166 AOI21X1_9/B 0 2.33fF
C167 AOI21X1_9/A 0 2.59fF
C168 NOR3X1_3/Y 0 2.04fF
C169 AOI22X1_6/B 0 2.56fF
C170 NAND3X1_59/Y 0 2.15fF
C171 OAI21X1_72/Y 0 2.33fF
C172 NAND3X1_62/Y 0 2.96fF
C173 NAND3X1_74/Y 0 2.18fF
C174 AOI22X1_11/A 0 2.12fF
C175 INVX1_39/Y 0 2.21fF
C176 AOI21X1_4/B 0 2.58fF
C177 OAI21X1_48/Y 0 2.14fF
C178 BUFX4_4/A 0 2.70fF
C179 INVX1_8/A 0 2.55fF
C180 AOI22X1_4/D 0 2.29fF
C181 NAND3X1_46/Y 0 2.23fF
C182 OAI21X1_43/C 0 2.13fF
C183 AOI22X1_6/D 0 3.02fF
C184 AOI22X1_6/C 0 2.23fF
C185 NAND2X1_79/Y 0 2.27fF
C186 NOR3X1_7/A 0 2.23fF
C187 INVX2_8/Y 0 2.02fF
C188 INVX1_39/A 0 2.10fF
C189 INVX4_4/Y 0 2.08fF
C190 INVX1_50/A 0 2.00fF
C191 OAI21X1_104/Y 0 2.01fF
C192 NAND2X1_110/Y 0 2.13fF
C193 INVX2_2/Y 0 2.17fF
C194 INVX1_18/A 0 2.02fF
C195 NAND3X1_9/Y 0 2.17fF
C196 AOI21X1_30/Y 0 2.04fF
C197 XNOR2X1_7/Y 0 2.17fF
C198 XNOR2X1_6/Y 0 2.29fF
C199 NAND3X1_96/A 0 2.23fF
C200 AND2X2_17/A 0 2.04fF
C201 AND2X2_16/Y 0 2.58fF
C202 NAND2X1_45/Y 0 2.10fF
C203 NAND3X1_7/Y 0 2.01fF
C204 OAI21X1_30/B 0 2.44fF
C205 NAND3X1_44/Y 0 2.16fF
C206 XNOR2X1_6/A 0 2.83fF
C207 NOR3X1_5/A 0 2.42fF
C208 NOR3X1_9/B 0 2.01fF
C209 OAI21X1_93/Y 0 2.58fF
C210 NAND3X1_89/Y 0 2.05fF
C211 NOR3X1_2/A 0 2.39fF
C212 NOR3X1_2/C 0 2.32fF
C213 INVX1_56/A 0 2.32fF
C214 INVX4_3/Y 0 2.36fF
C215 NAND2X1_39/Y 0 2.01fF
C216 NAND2X1_38/Y 0 2.18fF
C217 NAND3X1_32/Y 0 2.22fF
C218 INVX1_12/Y 0 2.10fF
C219 OAI22X1_5/B 0 2.78fF
C220 AND2X2_13/Y 0 2.04fF
C221 NAND3X1_90/Y 0 2.11fF
C222 NAND3X1_107/C 0 2.33fF
C223 AOI22X1_22/Y 0 2.03fF
C224 OAI21X1_122/Y 0 2.17fF
C225 OAI21X1_124/Y 0 2.06fF
C226 AND2X2_3/A 0 2.92fF
C227 NAND2X1_11/A 0 2.18fF
C228 OR2X2_2/B 0 3.04fF
C229 NAND3X1_6/Y 0 3.19fF
C230 OAI21X1_20/Y 0 2.00fF
C231 OAI22X1_5/A 0 2.06fF
C232 AOI21X1_44/A 0 2.09fF
C233 AOI22X1_14/D 0 2.41fF
C234 NAND2X1_119/A 0 2.02fF
C235 OAI22X1_6/Y 0 2.12fF
C236 NOR2X1_14/A 0 2.29fF
C237 OAI21X1_26/Y 0 2.31fF
C238 XOR2X1_2/A 0 2.00fF
C239 AOI22X1_9/D 0 2.27fF
C240 AOI21X1_82/B 0 2.68fF
C241 NOR3X1_1/B 0 2.26fF
C242 AOI21X1_72/B 0 3.00fF
C243 NOR2X1_4/B 0 2.22fF
C244 NAND3X1_2/Y 0 2.42fF
C245 OAI21X1_2/Y 0 2.41fF
C246 NOR2X1_9/A 0 2.23fF
C247 NAND3X1_22/B 0 2.38fF
C248 XNOR2X1_5/Y 0 2.34fF
C249 AOI21X1_70/B 0 2.12fF
C250 NOR2X1_6/Y 0 2.24fF
C251 INVX1_57/A 0 2.39fF
C252 NOR2X1_7/A 0 2.37fF
C253 AND2X2_5/B 0 2.09fF
C254 OR2X2_1/A 0 2.69fF
C255 AND2X2_5/Y 0 2.17fF
C256 NOR2X1_5/Y 0 2.11fF
C257 NAND3X1_3/B 0 2.28fF
C258 NAND3X1_1/Y 0 2.11fF
C259 NAND3X1_4/Y 0 2.17fF
