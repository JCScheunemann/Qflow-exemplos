module multiplicador (clk, A, B, S);

input clk;
input [7:0] A;
input [7:0] B;
output [15:0] S;

wire vdd = 1'b1;
wire gnd = 1'b0;

	BUFX4 BUFX4_1 ( .A(_85_), .Y(_85__bF_buf3) );
	BUFX4 BUFX4_2 ( .A(_85_), .Y(_85__bF_buf2) );
	BUFX4 BUFX4_3 ( .A(_85_), .Y(_85__bF_buf1) );
	BUFX4 BUFX4_4 ( .A(_85_), .Y(_85__bF_buf0) );
	NAND2X1 NAND2X1_1 ( .A(_276_), .B(_273_), .Y(_280_) );
	OAI21X1 OAI21X1_1 ( .A(_434_), .B(_275_), .C(_260_), .Y(_281_) );
	NAND3X1 NAND3X1_1 ( .A(_279_), .B(_280_), .C(_281_), .Y(_283_) );
	NAND2X1 NAND2X1_2 ( .A(_278_), .B(_283_), .Y(_284_) );
	NAND2X1 NAND2X1_3 ( .A(B[1]), .B(A[7]), .Y(_285_) );
	OAI22X1 OAI22X1_1 ( .A(_115_), .B(_285_), .C(_188_), .D(_193_), .Y(_286_) );
	AND2X2 AND2X2_1 ( .A(B[2]), .B(A[7]), .Y(_287_) );
	AOI22X1 AOI22X1_1 ( .A(B[1]), .B(A[7]), .C(B[2]), .D(A[6]), .Y(_288_) );
	AOI21X1 AOI21X1_1 ( .A(_108_), .B(_287_), .C(_288_), .Y(_289_) );
	NAND2X1 NAND2X1_4 ( .A(_289_), .B(_286_), .Y(_290_) );
	OR2X2 OR2X2_1 ( .A(_286_), .B(_289_), .Y(_291_) );
	NAND3X1 NAND3X1_2 ( .A(_290_), .B(_291_), .C(_284_), .Y(_292_) );
	NAND3X1 NAND3X1_3 ( .A(_279_), .B(_277_), .C(_274_), .Y(_294_) );
	NAND3X1 NAND3X1_4 ( .A(_272_), .B(_280_), .C(_281_), .Y(_295_) );
	NAND2X1 NAND2X1_5 ( .A(_294_), .B(_295_), .Y(_296_) );
	AND2X2 AND2X2_2 ( .A(_286_), .B(_289_), .Y(_297_) );
	NOR2X1 NOR2X1_1 ( .A(_289_), .B(_286_), .Y(_298_) );
	OAI21X1 OAI21X1_2 ( .A(_298_), .B(_297_), .C(_296_), .Y(_299_) );
	NAND2X1 NAND2X1_6 ( .A(_299_), .B(_292_), .Y(_300_) );
	NAND2X1 NAND2X1_7 ( .A(_269_), .B(_300_), .Y(_301_) );
	NOR3X1 NOR3X1_1 ( .A(_202_), .B(_203_), .C(_204_), .Y(_302_) );
	AOI21X1 AOI21X1_2 ( .A(_185_), .B(_205_), .C(_302_), .Y(_303_) );
	NAND3X1 NAND3X1_5 ( .A(_292_), .B(_299_), .C(_303_), .Y(_305_) );
	AOI22X1 AOI22X1_2 ( .A(_263_), .B(_267_), .C(_301_), .D(_305_), .Y(_306_) );
	NAND2X1 NAND2X1_8 ( .A(_263_), .B(_267_), .Y(_307_) );
	NAND3X1 NAND3X1_6 ( .A(_292_), .B(_299_), .C(_269_), .Y(_308_) );
	NAND2X1 NAND2X1_9 ( .A(_303_), .B(_300_), .Y(_309_) );
	AOI21X1 AOI21X1_3 ( .A(_309_), .B(_308_), .C(_307_), .Y(_310_) );
	OAI21X1 OAI21X1_3 ( .A(_310_), .B(_306_), .C(_254_), .Y(_311_) );
	NOR3X1 NOR3X1_2 ( .A(_216_), .B(_217_), .C(_215_), .Y(_312_) );
	AOI21X1 AOI21X1_4 ( .A(_173_), .B(_218_), .C(_312_), .Y(_313_) );
	NAND3X1 NAND3X1_7 ( .A(_307_), .B(_308_), .C(_309_), .Y(_314_) );
	AND2X2 AND2X2_3 ( .A(_267_), .B(_263_), .Y(_316_) );
	NAND3X1 NAND3X1_8 ( .A(_316_), .B(_301_), .C(_305_), .Y(_317_) );
	NAND3X1 NAND3X1_9 ( .A(_314_), .B(_317_), .C(_313_), .Y(_318_) );
	AOI21X1 AOI21X1_5 ( .A(_318_), .B(_311_), .C(_252_), .Y(_319_) );
	NAND3X1 NAND3X1_10 ( .A(_314_), .B(_317_), .C(_254_), .Y(_320_) );
	OAI21X1 OAI21X1_4 ( .A(_306_), .B(_310_), .C(_313_), .Y(_321_) );
	AOI21X1 AOI21X1_6 ( .A(_321_), .B(_320_), .C(_251_), .Y(_322_) );
	OAI21X1 OAI21X1_5 ( .A(_322_), .B(_319_), .C(_250_), .Y(_323_) );
	INVX1 INVX1_1 ( .A(_226_), .Y(_324_) );
	AOI21X1 AOI21X1_7 ( .A(_156_), .B(_232_), .C(_324_), .Y(_325_) );
	NAND3X1 NAND3X1_11 ( .A(_251_), .B(_320_), .C(_321_), .Y(_327_) );
	NAND3X1 NAND3X1_12 ( .A(_252_), .B(_311_), .C(_318_), .Y(_328_) );
	NAND3X1 NAND3X1_13 ( .A(_327_), .B(_328_), .C(_325_), .Y(_329_) );
	NAND2X1 NAND2X1_10 ( .A(_323_), .B(_329_), .Y(_330_) );
	XOR2X1 XOR2X1_1 ( .A(_246_), .B(_330_), .Y(_0__8_) );
	INVX1 INVX1_2 ( .A(_237_), .Y(_331_) );
	AOI21X1 AOI21X1_8 ( .A(_153_), .B(_240_), .C(_331_), .Y(_332_) );
	NAND3X1 NAND3X1_14 ( .A(_327_), .B(_328_), .C(_250_), .Y(_333_) );
	AOI21X1 AOI21X1_9 ( .A(_327_), .B(_328_), .C(_325_), .Y(_334_) );
	NOR3X1 NOR3X1_3 ( .A(_250_), .B(_322_), .C(_319_), .Y(_335_) );
	NOR2X1 NOR2X1_2 ( .A(_334_), .B(_335_), .Y(_337_) );
	OAI21X1 OAI21X1_6 ( .A(_337_), .B(_332_), .C(_333_), .Y(_338_) );
	AOI21X1 AOI21X1_10 ( .A(_317_), .B(_314_), .C(_254_), .Y(_339_) );
	OAI21X1 OAI21X1_7 ( .A(_252_), .B(_339_), .C(_320_), .Y(_340_) );
	NAND2X1 NAND2X1_11 ( .A(_262_), .B(_259_), .Y(_341_) );
	OAI21X1 OAI21X1_8 ( .A(_255_), .B(_341_), .C(_259_), .Y(_342_) );
	AOI21X1 AOI21X1_11 ( .A(_292_), .B(_299_), .C(_269_), .Y(_343_) );
	OAI21X1 OAI21X1_9 ( .A(_343_), .B(_316_), .C(_308_), .Y(_344_) );
	NAND2X1 NAND2X1_12 ( .A(A[2]), .B(B[7]), .Y(_345_) );
	NOR2X1 NOR2X1_3 ( .A(_521_), .B(_85__bF_buf3), .Y(_346_) );
	NOR2X1 NOR2X1_4 ( .A(_260_), .B(_273_), .Y(_347_) );
	OAI21X1 OAI21X1_10 ( .A(_272_), .B(_347_), .C(_274_), .Y(_348_) );
	NAND2X1 NAND2X1_13 ( .A(_346_), .B(_348_), .Y(_349_) );
	NAND2X1 NAND2X1_14 ( .A(B[3]), .B(A[5]), .Y(_350_) );
	NOR2X1 NOR2X1_5 ( .A(_276_), .B(_350_), .Y(_351_) );
	AOI21X1 AOI21X1_12 ( .A(_277_), .B(_279_), .C(_351_), .Y(_352_) );
	OAI21X1 OAI21X1_11 ( .A(_521_), .B(_85__bF_buf2), .C(_352_), .Y(_353_) );
	NAND3X1 NAND3X1_15 ( .A(_345_), .B(_353_), .C(_349_), .Y(_354_) );
	INVX1 INVX1_3 ( .A(_345_), .Y(_355_) );
	OAI21X1 OAI21X1_12 ( .A(_521_), .B(_85__bF_buf1), .C(_348_), .Y(_356_) );
	NAND2X1 NAND2X1_15 ( .A(_346_), .B(_352_), .Y(_358_) );
	NAND3X1 NAND3X1_16 ( .A(_355_), .B(_358_), .C(_356_), .Y(_359_) );
	NAND2X1 NAND2X1_16 ( .A(_354_), .B(_359_), .Y(_360_) );
	OAI21X1 OAI21X1_13 ( .A(_298_), .B(_296_), .C(_290_), .Y(_361_) );
	OAI21X1 OAI21X1_14 ( .A(_271_), .B(_110_), .C(_287_), .Y(_362_) );
	INVX1 INVX1_4 ( .A(_362_), .Y(_363_) );
	NAND2X1 NAND2X1_17 ( .A(A[4]), .B(B[5]), .Y(_364_) );
	INVX1 INVX1_5 ( .A(_364_), .Y(_365_) );
	AND2X2 AND2X2_4 ( .A(B[4]), .B(A[6]), .Y(_366_) );
	NAND2X1 NAND2X1_18 ( .A(_273_), .B(_366_), .Y(_367_) );
	NAND2X1 NAND2X1_19 ( .A(B[3]), .B(A[6]), .Y(_370_) );
	OAI21X1 OAI21X1_15 ( .A(_633_), .B(_275_), .C(_370_), .Y(_371_) );
	NAND3X1 NAND3X1_17 ( .A(_365_), .B(_371_), .C(_367_), .Y(_372_) );
	NAND2X1 NAND2X1_20 ( .A(B[4]), .B(A[6]), .Y(_373_) );
	NOR2X1 NOR2X1_6 ( .A(_350_), .B(_373_), .Y(_374_) );
	AOI22X1 AOI22X1_3 ( .A(B[3]), .B(A[6]), .C(B[4]), .D(A[5]), .Y(_375_) );
	OAI21X1 OAI21X1_16 ( .A(_375_), .B(_374_), .C(_364_), .Y(_376_) );
	NAND3X1 NAND3X1_18 ( .A(_363_), .B(_372_), .C(_376_), .Y(_377_) );
	NAND3X1 NAND3X1_19 ( .A(_364_), .B(_371_), .C(_367_), .Y(_378_) );
	OAI21X1 OAI21X1_17 ( .A(_375_), .B(_374_), .C(_365_), .Y(_379_) );
	NAND3X1 NAND3X1_20 ( .A(_362_), .B(_378_), .C(_379_), .Y(_381_) );
	AND2X2 AND2X2_5 ( .A(_377_), .B(_381_), .Y(_382_) );
	NAND2X1 NAND2X1_21 ( .A(_361_), .B(_382_), .Y(_383_) );
	AOI21X1 AOI21X1_13 ( .A(_284_), .B(_291_), .C(_297_), .Y(_384_) );
	NAND2X1 NAND2X1_22 ( .A(_377_), .B(_381_), .Y(_385_) );
	NAND2X1 NAND2X1_23 ( .A(_385_), .B(_384_), .Y(_386_) );
	NAND3X1 NAND3X1_21 ( .A(_386_), .B(_383_), .C(_360_), .Y(_387_) );
	NAND3X1 NAND3X1_22 ( .A(_355_), .B(_353_), .C(_349_), .Y(_388_) );
	NAND3X1 NAND3X1_23 ( .A(_345_), .B(_358_), .C(_356_), .Y(_389_) );
	NAND2X1 NAND2X1_24 ( .A(_388_), .B(_389_), .Y(_390_) );
	NOR2X1 NOR2X1_7 ( .A(_385_), .B(_384_), .Y(_392_) );
	NOR2X1 NOR2X1_8 ( .A(_361_), .B(_382_), .Y(_393_) );
	OAI21X1 OAI21X1_18 ( .A(_392_), .B(_393_), .C(_390_), .Y(_394_) );
	NAND3X1 NAND3X1_24 ( .A(_387_), .B(_394_), .C(_344_), .Y(_395_) );
	NOR2X1 NOR2X1_9 ( .A(_303_), .B(_300_), .Y(_396_) );
	AOI21X1 AOI21X1_14 ( .A(_307_), .B(_309_), .C(_396_), .Y(_397_) );
	NAND2X1 NAND2X1_25 ( .A(_385_), .B(_361_), .Y(_398_) );
	NAND2X1 NAND2X1_26 ( .A(_384_), .B(_382_), .Y(_399_) );
	AOI21X1 AOI21X1_15 ( .A(_399_), .B(_398_), .C(_390_), .Y(_400_) );
	AOI21X1 AOI21X1_16 ( .A(_383_), .B(_386_), .C(_360_), .Y(_401_) );
	OAI21X1 OAI21X1_19 ( .A(_401_), .B(_400_), .C(_397_), .Y(_403_) );
	NAND3X1 NAND3X1_25 ( .A(_342_), .B(_395_), .C(_403_), .Y(_404_) );
	INVX1 INVX1_6 ( .A(_342_), .Y(_405_) );
	OAI21X1 OAI21X1_20 ( .A(_401_), .B(_400_), .C(_344_), .Y(_406_) );
	NAND3X1 NAND3X1_26 ( .A(_387_), .B(_394_), .C(_397_), .Y(_407_) );
	NAND3X1 NAND3X1_27 ( .A(_405_), .B(_406_), .C(_407_), .Y(_408_) );
	NAND3X1 NAND3X1_28 ( .A(_404_), .B(_408_), .C(_340_), .Y(_409_) );
	AOI21X1 AOI21X1_17 ( .A(_408_), .B(_404_), .C(_340_), .Y(_410_) );
	INVX1 INVX1_7 ( .A(_410_), .Y(_411_) );
	NAND2X1 NAND2X1_27 ( .A(_409_), .B(_411_), .Y(_412_) );
	XNOR2X1 XNOR2X1_1 ( .A(_338_), .B(_412_), .Y(_0__9_) );
	AOI21X1 AOI21X1_18 ( .A(_407_), .B(_406_), .C(_405_), .Y(_414_) );
	AOI21X1 AOI21X1_19 ( .A(_403_), .B(_395_), .C(_342_), .Y(_415_) );
	OAI21X1 OAI21X1_21 ( .A(_415_), .B(_414_), .C(_340_), .Y(_416_) );
	INVX1 INVX1_8 ( .A(_320_), .Y(_417_) );
	AOI21X1 AOI21X1_20 ( .A(_251_), .B(_321_), .C(_417_), .Y(_418_) );
	NAND3X1 NAND3X1_29 ( .A(_404_), .B(_408_), .C(_418_), .Y(_419_) );
	AOI22X1 AOI22X1_4 ( .A(_419_), .B(_416_), .C(_323_), .D(_329_), .Y(_420_) );
	OAI21X1 OAI21X1_22 ( .A(_410_), .B(_333_), .C(_409_), .Y(_421_) );
	AOI21X1 AOI21X1_21 ( .A(_420_), .B(_246_), .C(_421_), .Y(_422_) );
	INVX1 INVX1_9 ( .A(_395_), .Y(_424_) );
	NAND2X1 NAND2X1_28 ( .A(_349_), .B(_388_), .Y(_425_) );
	OAI21X1 OAI21X1_23 ( .A(_390_), .B(_393_), .C(_383_), .Y(_426_) );
	NAND2X1 NAND2X1_29 ( .A(A[3]), .B(B[7]), .Y(_427_) );
	NOR2X1 NOR2X1_10 ( .A(_645_), .B(_85__bF_buf0), .Y(_428_) );
	OAI21X1 OAI21X1_24 ( .A(_364_), .B(_375_), .C(_367_), .Y(_429_) );
	NAND2X1 NAND2X1_30 ( .A(_428_), .B(_429_), .Y(_430_) );
	AOI22X1 AOI22X1_5 ( .A(_273_), .B(_366_), .C(_365_), .D(_371_), .Y(_431_) );
	OAI21X1 OAI21X1_25 ( .A(_645_), .B(_85__bF_buf3), .C(_431_), .Y(_432_) );
	NAND3X1 NAND3X1_30 ( .A(_427_), .B(_430_), .C(_432_), .Y(_433_) );
	INVX1 INVX1_10 ( .A(_427_), .Y(_435_) );
	NAND2X1 NAND2X1_31 ( .A(_430_), .B(_432_), .Y(_436_) );
	NAND2X1 NAND2X1_32 ( .A(_435_), .B(_436_), .Y(_437_) );
	NAND2X1 NAND2X1_33 ( .A(_433_), .B(_437_), .Y(_438_) );
	NAND2X1 NAND2X1_34 ( .A(_108_), .B(_287_), .Y(_439_) );
	NAND2X1 NAND2X1_35 ( .A(_439_), .B(_377_), .Y(_440_) );
	INVX2 INVX2_1 ( .A(B[5]), .Y(_441_) );
	NOR2X1 NOR2X1_11 ( .A(_275_), .B(_441_), .Y(_442_) );
	NAND2X1 NAND2X1_36 ( .A(B[4]), .B(A[7]), .Y(_443_) );
	INVX2 INVX2_2 ( .A(A[7]), .Y(_444_) );
	OAI21X1 OAI21X1_26 ( .A(_434_), .B(_444_), .C(_373_), .Y(_446_) );
	OAI21X1 OAI21X1_27 ( .A(_370_), .B(_443_), .C(_446_), .Y(_447_) );
	XOR2X1 XOR2X1_2 ( .A(_447_), .B(_442_), .Y(_448_) );
	INVX1 INVX1_11 ( .A(_448_), .Y(_449_) );
	NAND2X1 NAND2X1_37 ( .A(_440_), .B(_449_), .Y(_450_) );
	NAND3X1 NAND3X1_31 ( .A(_439_), .B(_377_), .C(_448_), .Y(_451_) );
	NAND3X1 NAND3X1_32 ( .A(_450_), .B(_451_), .C(_438_), .Y(_452_) );
	NAND3X1 NAND3X1_33 ( .A(_435_), .B(_430_), .C(_432_), .Y(_453_) );
	INVX2 INVX2_3 ( .A(B[7]), .Y(_454_) );
	OAI21X1 OAI21X1_28 ( .A(_521_), .B(_454_), .C(_436_), .Y(_455_) );
	NAND2X1 NAND2X1_38 ( .A(_453_), .B(_455_), .Y(_457_) );
	NAND2X1 NAND2X1_39 ( .A(_448_), .B(_440_), .Y(_458_) );
	OR2X2 OR2X2_2 ( .A(_440_), .B(_448_), .Y(_459_) );
	NAND3X1 NAND3X1_34 ( .A(_458_), .B(_459_), .C(_457_), .Y(_460_) );
	NAND3X1 NAND3X1_35 ( .A(_452_), .B(_460_), .C(_426_), .Y(_461_) );
	AOI21X1 AOI21X1_22 ( .A(_360_), .B(_386_), .C(_392_), .Y(_462_) );
	AOI21X1 AOI21X1_23 ( .A(_459_), .B(_458_), .C(_457_), .Y(_463_) );
	AOI21X1 AOI21X1_24 ( .A(_450_), .B(_451_), .C(_438_), .Y(_464_) );
	OAI21X1 OAI21X1_29 ( .A(_464_), .B(_463_), .C(_462_), .Y(_465_) );
	NAND3X1 NAND3X1_36 ( .A(_425_), .B(_461_), .C(_465_), .Y(_466_) );
	INVX1 INVX1_12 ( .A(_425_), .Y(_468_) );
	OAI21X1 OAI21X1_30 ( .A(_464_), .B(_463_), .C(_426_), .Y(_469_) );
	NAND3X1 NAND3X1_37 ( .A(_452_), .B(_462_), .C(_460_), .Y(_470_) );
	NAND3X1 NAND3X1_38 ( .A(_468_), .B(_470_), .C(_469_), .Y(_471_) );
	NAND2X1 NAND2X1_40 ( .A(_466_), .B(_471_), .Y(_472_) );
	OAI21X1 OAI21X1_31 ( .A(_424_), .B(_414_), .C(_472_), .Y(_473_) );
	AOI21X1 AOI21X1_25 ( .A(_342_), .B(_403_), .C(_424_), .Y(_474_) );
	NAND3X1 NAND3X1_39 ( .A(_466_), .B(_471_), .C(_474_), .Y(_475_) );
	NAND2X1 NAND2X1_41 ( .A(_475_), .B(_473_), .Y(_476_) );
	XNOR2X1 XNOR2X1_2 ( .A(_422_), .B(_476_), .Y(_0__10_) );
	NOR2X1 NOR2X1_12 ( .A(_474_), .B(_472_), .Y(_478_) );
	INVX1 INVX1_13 ( .A(_478_), .Y(_479_) );
	INVX1 INVX1_14 ( .A(_476_), .Y(_480_) );
	OAI21X1 OAI21X1_32 ( .A(_480_), .B(_422_), .C(_479_), .Y(_481_) );
	AOI21X1 AOI21X1_26 ( .A(_460_), .B(_452_), .C(_426_), .Y(_482_) );
	OAI21X1 OAI21X1_33 ( .A(_468_), .B(_482_), .C(_461_), .Y(_483_) );
	OAI21X1 OAI21X1_34 ( .A(_427_), .B(_436_), .C(_430_), .Y(_484_) );
	INVX1 INVX1_15 ( .A(_484_), .Y(_485_) );
	INVX1 INVX1_16 ( .A(_450_), .Y(_486_) );
	NOR2X1 NOR2X1_13 ( .A(_645_), .B(_454_), .Y(_487_) );
	INVX1 INVX1_17 ( .A(_487_), .Y(_488_) );
	NOR2X1 NOR2X1_14 ( .A(_370_), .B(_443_), .Y(_489_) );
	AOI21X1 AOI21X1_27 ( .A(_446_), .B(_442_), .C(_489_), .Y(_490_) );
	INVX1 INVX1_18 ( .A(_490_), .Y(_491_) );
	OAI21X1 OAI21X1_35 ( .A(_275_), .B(_85__bF_buf2), .C(_491_), .Y(_492_) );
	NAND2X1 NAND2X1_42 ( .A(A[5]), .B(B[6]), .Y(_493_) );
	INVX1 INVX1_19 ( .A(_493_), .Y(_494_) );
	NAND2X1 NAND2X1_43 ( .A(_494_), .B(_490_), .Y(_495_) );
	AOI21X1 AOI21X1_28 ( .A(_492_), .B(_495_), .C(_488_), .Y(_496_) );
	NAND2X1 NAND2X1_44 ( .A(_494_), .B(_491_), .Y(_497_) );
	OAI21X1 OAI21X1_36 ( .A(_275_), .B(_85__bF_buf1), .C(_490_), .Y(_500_) );
	AOI21X1 AOI21X1_29 ( .A(_497_), .B(_500_), .C(_487_), .Y(_501_) );
	NOR2X1 NOR2X1_15 ( .A(_441_), .B(_444_), .Y(_502_) );
	NAND2X1 NAND2X1_45 ( .A(_366_), .B(_502_), .Y(_503_) );
	OAI21X1 OAI21X1_37 ( .A(_441_), .B(_110_), .C(_443_), .Y(_504_) );
	NAND2X1 NAND2X1_46 ( .A(_504_), .B(_503_), .Y(_505_) );
	OAI21X1 OAI21X1_38 ( .A(_501_), .B(_496_), .C(_505_), .Y(_506_) );
	NAND3X1 NAND3X1_40 ( .A(_487_), .B(_500_), .C(_497_), .Y(_507_) );
	NAND3X1 NAND3X1_41 ( .A(_488_), .B(_495_), .C(_492_), .Y(_508_) );
	INVX1 INVX1_20 ( .A(_505_), .Y(_509_) );
	NAND3X1 NAND3X1_42 ( .A(_509_), .B(_507_), .C(_508_), .Y(_511_) );
	NAND2X1 NAND2X1_47 ( .A(_511_), .B(_506_), .Y(_512_) );
	OAI21X1 OAI21X1_39 ( .A(_486_), .B(_463_), .C(_512_), .Y(_513_) );
	AOI21X1 AOI21X1_30 ( .A(_438_), .B(_451_), .C(_486_), .Y(_514_) );
	NAND3X1 NAND3X1_43 ( .A(_506_), .B(_511_), .C(_514_), .Y(_515_) );
	AOI21X1 AOI21X1_31 ( .A(_515_), .B(_513_), .C(_485_), .Y(_516_) );
	INVX1 INVX1_21 ( .A(_451_), .Y(_517_) );
	OAI21X1 OAI21X1_40 ( .A(_517_), .B(_457_), .C(_450_), .Y(_518_) );
	NAND3X1 NAND3X1_44 ( .A(_506_), .B(_511_), .C(_518_), .Y(_519_) );
	NAND2X1 NAND2X1_48 ( .A(_512_), .B(_514_), .Y(_520_) );
	AOI21X1 AOI21X1_32 ( .A(_520_), .B(_519_), .C(_484_), .Y(_522_) );
	OAI21X1 OAI21X1_41 ( .A(_522_), .B(_516_), .C(_483_), .Y(_523_) );
	INVX1 INVX1_22 ( .A(_461_), .Y(_524_) );
	AOI21X1 AOI21X1_33 ( .A(_425_), .B(_465_), .C(_524_), .Y(_525_) );
	NAND3X1 NAND3X1_45 ( .A(_484_), .B(_519_), .C(_520_), .Y(_526_) );
	NAND3X1 NAND3X1_46 ( .A(_485_), .B(_513_), .C(_515_), .Y(_527_) );
	NAND3X1 NAND3X1_47 ( .A(_526_), .B(_527_), .C(_525_), .Y(_528_) );
	NAND3X1 NAND3X1_48 ( .A(_523_), .B(_528_), .C(_481_), .Y(_529_) );
	AND2X2 AND2X2_6 ( .A(_420_), .B(_246_), .Y(_530_) );
	OAI21X1 OAI21X1_42 ( .A(_421_), .B(_530_), .C(_476_), .Y(_531_) );
	NAND2X1 NAND2X1_49 ( .A(_528_), .B(_523_), .Y(_533_) );
	NAND3X1 NAND3X1_49 ( .A(_479_), .B(_533_), .C(_531_), .Y(_534_) );
	NAND2X1 NAND2X1_50 ( .A(_534_), .B(_529_), .Y(_0__11_) );
	OAI21X1 OAI21X1_43 ( .A(_514_), .B(_512_), .C(_526_), .Y(_535_) );
	OAI21X1 OAI21X1_44 ( .A(_493_), .B(_490_), .C(_507_), .Y(_536_) );
	OAI21X1 OAI21X1_45 ( .A(_110_), .B(_85__bF_buf0), .C(_503_), .Y(_537_) );
	OAI21X1 OAI21X1_46 ( .A(_85__bF_buf3), .B(_503_), .C(_537_), .Y(_538_) );
	OAI21X1 OAI21X1_47 ( .A(_275_), .B(_454_), .C(_538_), .Y(_539_) );
	NAND2X1 NAND2X1_51 ( .A(A[5]), .B(B[7]), .Y(_540_) );
	OR2X2 OR2X2_3 ( .A(_538_), .B(_540_), .Y(_541_) );
	NAND3X1 NAND3X1_50 ( .A(_502_), .B(_539_), .C(_541_), .Y(_543_) );
	NAND2X1 NAND2X1_52 ( .A(_539_), .B(_541_), .Y(_544_) );
	OAI21X1 OAI21X1_48 ( .A(_441_), .B(_444_), .C(_544_), .Y(_545_) );
	NAND2X1 NAND2X1_53 ( .A(_543_), .B(_545_), .Y(_546_) );
	OR2X2 OR2X2_4 ( .A(_546_), .B(_511_), .Y(_547_) );
	NAND2X1 NAND2X1_54 ( .A(_511_), .B(_546_), .Y(_548_) );
	NAND3X1 NAND3X1_51 ( .A(_536_), .B(_548_), .C(_547_), .Y(_549_) );
	INVX1 INVX1_23 ( .A(_536_), .Y(_550_) );
	NOR2X1 NOR2X1_16 ( .A(_511_), .B(_546_), .Y(_551_) );
	AND2X2 AND2X2_7 ( .A(_546_), .B(_511_), .Y(_552_) );
	OAI21X1 OAI21X1_49 ( .A(_551_), .B(_552_), .C(_550_), .Y(_554_) );
	AOI21X1 AOI21X1_34 ( .A(_554_), .B(_549_), .C(_535_), .Y(_555_) );
	INVX1 INVX1_24 ( .A(_555_), .Y(_556_) );
	INVX1 INVX1_25 ( .A(_535_), .Y(_557_) );
	NAND2X1 NAND2X1_55 ( .A(_549_), .B(_554_), .Y(_558_) );
	OR2X2 OR2X2_5 ( .A(_558_), .B(_557_), .Y(_559_) );
	NAND2X1 NAND2X1_56 ( .A(_556_), .B(_559_), .Y(_560_) );
	OAI21X1 OAI21X1_50 ( .A(_522_), .B(_516_), .C(_525_), .Y(_561_) );
	NAND2X1 NAND2X1_57 ( .A(_526_), .B(_527_), .Y(_562_) );
	OAI22X1 OAI22X1_2 ( .A(_474_), .B(_472_), .C(_525_), .D(_562_), .Y(_563_) );
	AOI22X1 AOI22X1_6 ( .A(_523_), .B(_528_), .C(_473_), .D(_475_), .Y(_565_) );
	AOI22X1 AOI22X1_7 ( .A(_561_), .B(_563_), .C(_421_), .D(_565_), .Y(_566_) );
	NAND3X1 NAND3X1_52 ( .A(_565_), .B(_246_), .C(_420_), .Y(_567_) );
	AOI21X1 AOI21X1_35 ( .A(_567_), .B(_566_), .C(_560_), .Y(_568_) );
	NOR2X1 NOR2X1_17 ( .A(_557_), .B(_558_), .Y(_569_) );
	NOR2X1 NOR2X1_18 ( .A(_555_), .B(_569_), .Y(_570_) );
	NAND2X1 NAND2X1_58 ( .A(_561_), .B(_563_), .Y(_571_) );
	NAND2X1 NAND2X1_59 ( .A(_533_), .B(_476_), .Y(_572_) );
	NAND2X1 NAND2X1_60 ( .A(_571_), .B(_572_), .Y(_573_) );
	AOI21X1 AOI21X1_36 ( .A(_404_), .B(_408_), .C(_418_), .Y(_574_) );
	NAND2X1 NAND2X1_61 ( .A(_404_), .B(_408_), .Y(_576_) );
	NOR2X1 NOR2X1_19 ( .A(_340_), .B(_576_), .Y(_577_) );
	OAI22X1 OAI22X1_3 ( .A(_574_), .B(_577_), .C(_334_), .D(_335_), .Y(_578_) );
	OAI21X1 OAI21X1_51 ( .A(_418_), .B(_576_), .C(_333_), .Y(_579_) );
	AOI22X1 AOI22X1_8 ( .A(_563_), .B(_561_), .C(_411_), .D(_579_), .Y(_580_) );
	OAI21X1 OAI21X1_52 ( .A(_332_), .B(_578_), .C(_580_), .Y(_581_) );
	AOI21X1 AOI21X1_37 ( .A(_581_), .B(_573_), .C(_570_), .Y(_582_) );
	NOR2X1 NOR2X1_20 ( .A(_568_), .B(_582_), .Y(_0__12_) );
	NAND3X1 NAND3X1_53 ( .A(_570_), .B(_573_), .C(_581_), .Y(_583_) );
	OAI21X1 OAI21X1_53 ( .A(_550_), .B(_552_), .C(_547_), .Y(_584_) );
	OAI21X1 OAI21X1_54 ( .A(_85__bF_buf2), .B(_503_), .C(_541_), .Y(_586_) );
	NOR2X1 NOR2X1_21 ( .A(_110_), .B(_85__bF_buf1), .Y(_587_) );
	NOR2X1 NOR2X1_22 ( .A(_444_), .B(_454_), .Y(_588_) );
	NAND2X1 NAND2X1_62 ( .A(_587_), .B(_588_), .Y(_589_) );
	OAI22X1 OAI22X1_4 ( .A(_110_), .B(_454_), .C(_85__bF_buf0), .D(_444_), .Y(_590_) );
	NAND2X1 NAND2X1_63 ( .A(_590_), .B(_589_), .Y(_591_) );
	NAND2X1 NAND2X1_64 ( .A(_591_), .B(_543_), .Y(_592_) );
	OR2X2 OR2X2_6 ( .A(_543_), .B(_591_), .Y(_593_) );
	NAND2X1 NAND2X1_65 ( .A(_592_), .B(_593_), .Y(_594_) );
	XNOR2X1 XNOR2X1_3 ( .A(_594_), .B(_586_), .Y(_595_) );
	NAND2X1 NAND2X1_66 ( .A(_584_), .B(_595_), .Y(_597_) );
	AOI21X1 AOI21X1_38 ( .A(_536_), .B(_548_), .C(_551_), .Y(_598_) );
	XOR2X1 XOR2X1_3 ( .A(_594_), .B(_586_), .Y(_599_) );
	NAND2X1 NAND2X1_67 ( .A(_598_), .B(_599_), .Y(_600_) );
	AND2X2 AND2X2_8 ( .A(_600_), .B(_597_), .Y(_601_) );
	NAND3X1 NAND3X1_54 ( .A(_559_), .B(_601_), .C(_583_), .Y(_602_) );
	NAND2X1 NAND2X1_68 ( .A(_597_), .B(_600_), .Y(_603_) );
	OAI21X1 OAI21X1_55 ( .A(_569_), .B(_568_), .C(_603_), .Y(_604_) );
	NAND2X1 NAND2X1_69 ( .A(_604_), .B(_602_), .Y(_0__13_) );
	NOR3X1 NOR3X1_4 ( .A(_555_), .B(_603_), .C(_569_), .Y(_605_) );
	NAND3X1 NAND3X1_55 ( .A(_573_), .B(_605_), .C(_581_), .Y(_607_) );
	OAI21X1 OAI21X1_56 ( .A(_603_), .B(_559_), .C(_597_), .Y(_608_) );
	INVX1 INVX1_26 ( .A(_608_), .Y(_609_) );
	INVX1 INVX1_27 ( .A(_593_), .Y(_610_) );
	AOI21X1 AOI21X1_39 ( .A(_586_), .B(_592_), .C(_610_), .Y(_611_) );
	OAI21X1 OAI21X1_57 ( .A(_110_), .B(_85__bF_buf3), .C(_588_), .Y(_612_) );
	XOR2X1 XOR2X1_4 ( .A(_611_), .B(_612_), .Y(_613_) );
	NAND3X1 NAND3X1_56 ( .A(_609_), .B(_613_), .C(_607_), .Y(_614_) );
	NAND3X1 NAND3X1_57 ( .A(_556_), .B(_601_), .C(_559_), .Y(_615_) );
	AOI21X1 AOI21X1_40 ( .A(_567_), .B(_566_), .C(_615_), .Y(_616_) );
	INVX1 INVX1_28 ( .A(_613_), .Y(_618_) );
	OAI21X1 OAI21X1_58 ( .A(_608_), .B(_616_), .C(_618_), .Y(_619_) );
	NAND2X1 NAND2X1_70 ( .A(_619_), .B(_614_), .Y(_0__14_) );
	OAI21X1 OAI21X1_59 ( .A(_608_), .B(_616_), .C(_613_), .Y(_620_) );
	NOR2X1 NOR2X1_23 ( .A(_612_), .B(_611_), .Y(_621_) );
	AOI21X1 AOI21X1_41 ( .A(_587_), .B(_588_), .C(_621_), .Y(_622_) );
	NAND2X1 NAND2X1_71 ( .A(_622_), .B(_620_), .Y(_0__15_) );
	NOR2X1 NOR2X1_24 ( .A(_270_), .B(_228_), .Y(_0__0_) );
	INVX1 INVX1_29 ( .A(_293_), .Y(_623_) );
	NOR2X1 NOR2X1_25 ( .A(_249_), .B(_282_), .Y(_624_) );
	NOR2X1 NOR2X1_26 ( .A(_624_), .B(_623_), .Y(_0__1_) );
	XNOR2X1 XNOR2X1_4 ( .A(_402_), .B(_623_), .Y(_0__2_) );
	BUFX2 BUFX2_1 ( .A(_654__0_), .Y(S[0]) );
	BUFX2 BUFX2_2 ( .A(_654__1_), .Y(S[1]) );
	BUFX2 BUFX2_3 ( .A(_654__2_), .Y(S[2]) );
	BUFX2 BUFX2_4 ( .A(_654__3_), .Y(S[3]) );
	BUFX2 BUFX2_5 ( .A(_654__4_), .Y(S[4]) );
	BUFX2 BUFX2_6 ( .A(_654__5_), .Y(S[5]) );
	BUFX2 BUFX2_7 ( .A(_654__6_), .Y(S[6]) );
	BUFX2 BUFX2_8 ( .A(_654__7_), .Y(S[7]) );
	BUFX2 BUFX2_9 ( .A(_654__8_), .Y(S[8]) );
	BUFX2 BUFX2_10 ( .A(_654__9_), .Y(S[9]) );
	BUFX2 BUFX2_11 ( .A(_654__10_), .Y(S[10]) );
	BUFX2 BUFX2_12 ( .A(_654__11_), .Y(S[11]) );
	BUFX2 BUFX2_13 ( .A(_654__12_), .Y(S[12]) );
	BUFX2 BUFX2_14 ( .A(_654__13_), .Y(S[13]) );
	BUFX2 BUFX2_15 ( .A(_654__14_), .Y(S[14]) );
	BUFX2 BUFX2_16 ( .A(_654__15_), .Y(S[15]) );
	DFFPOSX1 DFFPOSX1_1 ( .CLK(clk), .D(_0__13_), .Q(_654__13_) );
	DFFPOSX1 DFFPOSX1_2 ( .CLK(clk), .D(_0__14_), .Q(_654__14_) );
	DFFPOSX1 DFFPOSX1_3 ( .CLK(clk), .D(_0__15_), .Q(_654__15_) );
	DFFPOSX1 DFFPOSX1_4 ( .CLK(clk), .D(_0__0_), .Q(_654__0_) );
	DFFPOSX1 DFFPOSX1_5 ( .CLK(clk), .D(_0__1_), .Q(_654__1_) );
	DFFPOSX1 DFFPOSX1_6 ( .CLK(clk), .D(_0__2_), .Q(_654__2_) );
	DFFPOSX1 DFFPOSX1_7 ( .CLK(clk), .D(_0__3_), .Q(_654__3_) );
	DFFPOSX1 DFFPOSX1_8 ( .CLK(clk), .D(_0__4_), .Q(_654__4_) );
	DFFPOSX1 DFFPOSX1_9 ( .CLK(clk), .D(_0__5_), .Q(_654__5_) );
	DFFPOSX1 DFFPOSX1_10 ( .CLK(clk), .D(_0__6_), .Q(_654__6_) );
	DFFPOSX1 DFFPOSX1_11 ( .CLK(clk), .D(_0__7_), .Q(_654__7_) );
	DFFPOSX1 DFFPOSX1_12 ( .CLK(clk), .D(_0__8_), .Q(_654__8_) );
	DFFPOSX1 DFFPOSX1_13 ( .CLK(clk), .D(_0__9_), .Q(_654__9_) );
	DFFPOSX1 DFFPOSX1_14 ( .CLK(clk), .D(_0__10_), .Q(_654__10_) );
	DFFPOSX1 DFFPOSX1_15 ( .CLK(clk), .D(_0__11_), .Q(_654__11_) );
	DFFPOSX1 DFFPOSX1_16 ( .CLK(clk), .D(_0__12_), .Q(_654__12_) );
	INVX2 INVX2_4 ( .A(B[0]), .Y(_228_) );
	INVX2 INVX2_5 ( .A(A[1]), .Y(_248_) );
	NOR2X1 NOR2X1_27 ( .A(_228_), .B(_248_), .Y(_249_) );
	INVX2 INVX2_6 ( .A(A[0]), .Y(_270_) );
	INVX2 INVX2_7 ( .A(B[1]), .Y(_271_) );
	NOR2X1 NOR2X1_28 ( .A(_270_), .B(_271_), .Y(_282_) );
	NAND2X1 NAND2X1_72 ( .A(_249_), .B(_282_), .Y(_293_) );
	INVX1 INVX1_30 ( .A(B[2]), .Y(_304_) );
	NOR2X1 NOR2X1_29 ( .A(_270_), .B(_304_), .Y(_315_) );
	INVX1 INVX1_31 ( .A(_315_), .Y(_326_) );
	NAND2X1 NAND2X1_73 ( .A(B[1]), .B(A[2]), .Y(_336_) );
	INVX1 INVX1_32 ( .A(_336_), .Y(_357_) );
	NAND2X1 NAND2X1_74 ( .A(_357_), .B(_249_), .Y(_368_) );
	NAND2X1 NAND2X1_75 ( .A(B[0]), .B(A[2]), .Y(_369_) );
	OAI21X1 OAI21X1_60 ( .A(_271_), .B(_248_), .C(_369_), .Y(_380_) );
	NAND2X1 NAND2X1_76 ( .A(_380_), .B(_368_), .Y(_391_) );
	XNOR2X1 XNOR2X1_5 ( .A(_391_), .B(_326_), .Y(_402_) );
	NOR2X1 NOR2X1_30 ( .A(_293_), .B(_402_), .Y(_413_) );
	INVX1 INVX1_33 ( .A(_413_), .Y(_423_) );
	INVX4 INVX4_1 ( .A(B[3]), .Y(_434_) );
	NOR2X1 NOR2X1_31 ( .A(_434_), .B(_270_), .Y(_445_) );
	INVX2 INVX2_8 ( .A(_445_), .Y(_456_) );
	AOI22X1 AOI22X1_9 ( .A(_249_), .B(_357_), .C(_315_), .D(_380_), .Y(_467_) );
	INVX1 INVX1_34 ( .A(_467_), .Y(_477_) );
	NAND2X1 NAND2X1_77 ( .A(B[2]), .B(A[1]), .Y(_498_) );
	INVX1 INVX1_35 ( .A(_498_), .Y(_499_) );
	NAND2X1 NAND2X1_78 ( .A(B[1]), .B(A[3]), .Y(_510_) );
	INVX4 INVX4_2 ( .A(A[3]), .Y(_521_) );
	OAI21X1 OAI21X1_61 ( .A(_228_), .B(_521_), .C(_336_), .Y(_532_) );
	OAI21X1 OAI21X1_62 ( .A(_369_), .B(_510_), .C(_532_), .Y(_542_) );
	XNOR2X1 XNOR2X1_6 ( .A(_542_), .B(_499_), .Y(_553_) );
	NAND2X1 NAND2X1_79 ( .A(_477_), .B(_553_), .Y(_564_) );
	XNOR2X1 XNOR2X1_7 ( .A(_542_), .B(_498_), .Y(_575_) );
	NAND2X1 NAND2X1_80 ( .A(_467_), .B(_575_), .Y(_585_) );
	NAND3X1 NAND3X1_58 ( .A(_456_), .B(_585_), .C(_564_), .Y(_596_) );
	NOR2X1 NOR2X1_32 ( .A(_467_), .B(_575_), .Y(_606_) );
	NOR2X1 NOR2X1_33 ( .A(_477_), .B(_553_), .Y(_617_) );
	OAI21X1 OAI21X1_63 ( .A(_606_), .B(_617_), .C(_445_), .Y(_625_) );
	AOI21X1 AOI21X1_42 ( .A(_625_), .B(_596_), .C(_423_), .Y(_626_) );
	NAND3X1 NAND3X1_59 ( .A(_445_), .B(_585_), .C(_564_), .Y(_627_) );
	OAI21X1 OAI21X1_64 ( .A(_606_), .B(_617_), .C(_456_), .Y(_628_) );
	AOI21X1 AOI21X1_43 ( .A(_628_), .B(_627_), .C(_413_), .Y(_629_) );
	NOR2X1 NOR2X1_34 ( .A(_626_), .B(_629_), .Y(_0__3_) );
	NAND3X1 NAND3X1_60 ( .A(_413_), .B(_627_), .C(_628_), .Y(_630_) );
	OAI21X1 OAI21X1_65 ( .A(_456_), .B(_617_), .C(_564_), .Y(_631_) );
	NAND2X1 NAND2X1_81 ( .A(A[1]), .B(B[4]), .Y(_632_) );
	INVX2 INVX2_9 ( .A(B[4]), .Y(_633_) );
	NAND2X1 NAND2X1_82 ( .A(B[3]), .B(A[1]), .Y(_634_) );
	OAI21X1 OAI21X1_66 ( .A(_270_), .B(_633_), .C(_634_), .Y(_635_) );
	OAI21X1 OAI21X1_67 ( .A(_632_), .B(_456_), .C(_635_), .Y(_636_) );
	NAND2X1 NAND2X1_83 ( .A(B[0]), .B(A[3]), .Y(_637_) );
	AND2X2 AND2X2_9 ( .A(_336_), .B(_637_), .Y(_638_) );
	OAI22X1 OAI22X1_5 ( .A(_369_), .B(_510_), .C(_498_), .D(_638_), .Y(_639_) );
	NAND2X1 NAND2X1_84 ( .A(B[2]), .B(A[2]), .Y(_640_) );
	INVX1 INVX1_36 ( .A(_640_), .Y(_641_) );
	AND2X2 AND2X2_10 ( .A(B[1]), .B(A[3]), .Y(_642_) );
	AND2X2 AND2X2_11 ( .A(A[4]), .B(B[0]), .Y(_643_) );
	NAND2X1 NAND2X1_85 ( .A(_642_), .B(_643_), .Y(_644_) );
	INVX4 INVX4_3 ( .A(A[4]), .Y(_645_) );
	OAI21X1 OAI21X1_68 ( .A(_645_), .B(_228_), .C(_510_), .Y(_646_) );
	NAND3X1 NAND3X1_61 ( .A(_641_), .B(_646_), .C(_644_), .Y(_647_) );
	NAND2X1 NAND2X1_86 ( .A(A[4]), .B(B[0]), .Y(_648_) );
	NOR2X1 NOR2X1_35 ( .A(_510_), .B(_648_), .Y(_649_) );
	AND2X2 AND2X2_12 ( .A(_510_), .B(_648_), .Y(_650_) );
	OAI21X1 OAI21X1_69 ( .A(_649_), .B(_650_), .C(_640_), .Y(_651_) );
	NAND3X1 NAND3X1_62 ( .A(_647_), .B(_651_), .C(_639_), .Y(_652_) );
	NOR2X1 NOR2X1_36 ( .A(_336_), .B(_637_), .Y(_653_) );
	AOI21X1 AOI21X1_44 ( .A(_532_), .B(_499_), .C(_653_), .Y(_1_) );
	OAI21X1 OAI21X1_70 ( .A(_271_), .B(_521_), .C(_643_), .Y(_2_) );
	OAI21X1 OAI21X1_71 ( .A(_645_), .B(_228_), .C(_642_), .Y(_3_) );
	AOI21X1 AOI21X1_45 ( .A(_2_), .B(_3_), .C(_640_), .Y(_4_) );
	AOI21X1 AOI21X1_46 ( .A(_644_), .B(_646_), .C(_641_), .Y(_5_) );
	OAI21X1 OAI21X1_72 ( .A(_5_), .B(_4_), .C(_1_), .Y(_6_) );
	NAND2X1 NAND2X1_87 ( .A(_652_), .B(_6_), .Y(_7_) );
	NOR2X1 NOR2X1_37 ( .A(_636_), .B(_7_), .Y(_8_) );
	INVX1 INVX1_37 ( .A(_636_), .Y(_9_) );
	AOI21X1 AOI21X1_47 ( .A(_6_), .B(_652_), .C(_9_), .Y(_10_) );
	OAI21X1 OAI21X1_73 ( .A(_8_), .B(_10_), .C(_631_), .Y(_11_) );
	AOI21X1 AOI21X1_48 ( .A(_585_), .B(_445_), .C(_606_), .Y(_12_) );
	OR2X2 OR2X2_7 ( .A(_7_), .B(_636_), .Y(_13_) );
	INVX1 INVX1_38 ( .A(_10_), .Y(_14_) );
	NAND3X1 NAND3X1_63 ( .A(_14_), .B(_13_), .C(_12_), .Y(_15_) );
	AOI21X1 AOI21X1_49 ( .A(_11_), .B(_15_), .C(_630_), .Y(_16_) );
	NAND3X1 NAND3X1_64 ( .A(_13_), .B(_14_), .C(_631_), .Y(_17_) );
	OAI21X1 OAI21X1_74 ( .A(_8_), .B(_10_), .C(_12_), .Y(_18_) );
	AOI21X1 AOI21X1_50 ( .A(_17_), .B(_18_), .C(_626_), .Y(_19_) );
	NOR2X1 NOR2X1_38 ( .A(_16_), .B(_19_), .Y(_0__4_) );
	NAND3X1 NAND3X1_65 ( .A(_18_), .B(_17_), .C(_626_), .Y(_20_) );
	INVX1 INVX1_39 ( .A(_632_), .Y(_21_) );
	NAND2X1 NAND2X1_88 ( .A(_21_), .B(_445_), .Y(_22_) );
	INVX1 INVX1_40 ( .A(_22_), .Y(_23_) );
	AOI21X1 AOI21X1_51 ( .A(_651_), .B(_647_), .C(_639_), .Y(_24_) );
	OAI21X1 OAI21X1_75 ( .A(_636_), .B(_24_), .C(_652_), .Y(_25_) );
	NAND2X1 NAND2X1_89 ( .A(A[0]), .B(B[5]), .Y(_26_) );
	INVX4 INVX4_4 ( .A(A[2]), .Y(_27_) );
	NOR2X1 NOR2X1_39 ( .A(_434_), .B(_27_), .Y(_28_) );
	NAND2X1 NAND2X1_90 ( .A(_21_), .B(_28_), .Y(_29_) );
	OAI21X1 OAI21X1_76 ( .A(_434_), .B(_27_), .C(_632_), .Y(_30_) );
	NAND3X1 NAND3X1_66 ( .A(_26_), .B(_30_), .C(_29_), .Y(_31_) );
	INVX1 INVX1_41 ( .A(_26_), .Y(_32_) );
	NAND2X1 NAND2X1_91 ( .A(A[2]), .B(B[4]), .Y(_33_) );
	OAI21X1 OAI21X1_77 ( .A(_634_), .B(_33_), .C(_30_), .Y(_34_) );
	NAND2X1 NAND2X1_92 ( .A(_32_), .B(_34_), .Y(_35_) );
	NAND2X1 NAND2X1_93 ( .A(_31_), .B(_35_), .Y(_36_) );
	OAI21X1 OAI21X1_78 ( .A(_640_), .B(_650_), .C(_644_), .Y(_37_) );
	NAND2X1 NAND2X1_94 ( .A(A[3]), .B(B[2]), .Y(_38_) );
	INVX1 INVX1_42 ( .A(_38_), .Y(_39_) );
	AND2X2 AND2X2_13 ( .A(A[4]), .B(B[1]), .Y(_40_) );
	AND2X2 AND2X2_14 ( .A(B[0]), .B(A[5]), .Y(_41_) );
	NAND2X1 NAND2X1_95 ( .A(_40_), .B(_41_), .Y(_42_) );
	NAND2X1 NAND2X1_96 ( .A(B[0]), .B(A[5]), .Y(_43_) );
	OAI21X1 OAI21X1_79 ( .A(_645_), .B(_271_), .C(_43_), .Y(_44_) );
	NAND3X1 NAND3X1_67 ( .A(_39_), .B(_44_), .C(_42_), .Y(_45_) );
	OAI21X1 OAI21X1_80 ( .A(_645_), .B(_271_), .C(_41_), .Y(_46_) );
	NAND2X1 NAND2X1_97 ( .A(_43_), .B(_40_), .Y(_47_) );
	NAND3X1 NAND3X1_68 ( .A(_38_), .B(_47_), .C(_46_), .Y(_48_) );
	NAND3X1 NAND3X1_69 ( .A(_45_), .B(_48_), .C(_37_), .Y(_49_) );
	AOI21X1 AOI21X1_52 ( .A(_646_), .B(_641_), .C(_649_), .Y(_50_) );
	AOI21X1 AOI21X1_53 ( .A(_46_), .B(_47_), .C(_38_), .Y(_51_) );
	AOI22X1 AOI22X1_10 ( .A(A[3]), .B(B[2]), .C(_44_), .D(_42_), .Y(_52_) );
	OAI21X1 OAI21X1_81 ( .A(_52_), .B(_51_), .C(_50_), .Y(_53_) );
	NAND3X1 NAND3X1_70 ( .A(_49_), .B(_53_), .C(_36_), .Y(_54_) );
	NAND3X1 NAND3X1_71 ( .A(_32_), .B(_30_), .C(_29_), .Y(_55_) );
	NAND3X1 NAND3X1_72 ( .A(B[3]), .B(A[2]), .C(_632_), .Y(_56_) );
	OAI21X1 OAI21X1_82 ( .A(_434_), .B(_27_), .C(_21_), .Y(_57_) );
	NAND3X1 NAND3X1_73 ( .A(_26_), .B(_56_), .C(_57_), .Y(_58_) );
	NAND2X1 NAND2X1_98 ( .A(_58_), .B(_55_), .Y(_59_) );
	OAI21X1 OAI21X1_83 ( .A(_52_), .B(_51_), .C(_37_), .Y(_60_) );
	NAND3X1 NAND3X1_74 ( .A(_45_), .B(_48_), .C(_50_), .Y(_61_) );
	NAND3X1 NAND3X1_75 ( .A(_61_), .B(_59_), .C(_60_), .Y(_62_) );
	NAND3X1 NAND3X1_76 ( .A(_62_), .B(_54_), .C(_25_), .Y(_63_) );
	NOR3X1 NOR3X1_5 ( .A(_1_), .B(_5_), .C(_4_), .Y(_64_) );
	AOI21X1 AOI21X1_54 ( .A(_9_), .B(_6_), .C(_64_), .Y(_65_) );
	AOI22X1 AOI22X1_11 ( .A(_31_), .B(_35_), .C(_61_), .D(_60_), .Y(_66_) );
	AOI21X1 AOI21X1_55 ( .A(_53_), .B(_49_), .C(_36_), .Y(_67_) );
	OAI21X1 OAI21X1_84 ( .A(_66_), .B(_67_), .C(_65_), .Y(_68_) );
	NAND3X1 NAND3X1_77 ( .A(_23_), .B(_63_), .C(_68_), .Y(_69_) );
	OAI21X1 OAI21X1_85 ( .A(_66_), .B(_67_), .C(_25_), .Y(_70_) );
	NAND3X1 NAND3X1_78 ( .A(_54_), .B(_62_), .C(_65_), .Y(_71_) );
	NAND3X1 NAND3X1_79 ( .A(_22_), .B(_71_), .C(_70_), .Y(_72_) );
	NAND3X1 NAND3X1_80 ( .A(_69_), .B(_17_), .C(_72_), .Y(_73_) );
	NOR3X1 NOR3X1_6 ( .A(_8_), .B(_10_), .C(_12_), .Y(_74_) );
	NAND3X1 NAND3X1_81 ( .A(_22_), .B(_63_), .C(_68_), .Y(_75_) );
	NAND3X1 NAND3X1_82 ( .A(_23_), .B(_71_), .C(_70_), .Y(_76_) );
	NAND3X1 NAND3X1_83 ( .A(_75_), .B(_76_), .C(_74_), .Y(_77_) );
	AOI21X1 AOI21X1_56 ( .A(_77_), .B(_73_), .C(_20_), .Y(_78_) );
	NAND3X1 NAND3X1_84 ( .A(_69_), .B(_72_), .C(_74_), .Y(_79_) );
	NAND3X1 NAND3X1_85 ( .A(_75_), .B(_17_), .C(_76_), .Y(_80_) );
	AOI21X1 AOI21X1_57 ( .A(_79_), .B(_80_), .C(_16_), .Y(_81_) );
	NOR2X1 NOR2X1_40 ( .A(_78_), .B(_81_), .Y(_0__5_) );
	AOI21X1 AOI21X1_58 ( .A(_76_), .B(_75_), .C(_17_), .Y(_82_) );
	AOI21X1 AOI21X1_59 ( .A(_54_), .B(_62_), .C(_25_), .Y(_83_) );
	OAI21X1 OAI21X1_86 ( .A(_22_), .B(_83_), .C(_63_), .Y(_84_) );
	INVX8 INVX8_1 ( .A(B[6]), .Y(_85_) );
	OAI21X1 OAI21X1_87 ( .A(_26_), .B(_34_), .C(_29_), .Y(_86_) );
	OAI21X1 OAI21X1_88 ( .A(_270_), .B(_85__bF_buf2), .C(_86_), .Y(_87_) );
	NOR2X1 NOR2X1_41 ( .A(_270_), .B(_85__bF_buf1), .Y(_88_) );
	NAND3X1 NAND3X1_86 ( .A(_29_), .B(_88_), .C(_55_), .Y(_89_) );
	NAND2X1 NAND2X1_99 ( .A(_89_), .B(_87_), .Y(_90_) );
	AOI21X1 AOI21X1_60 ( .A(_48_), .B(_45_), .C(_37_), .Y(_91_) );
	OAI21X1 OAI21X1_89 ( .A(_91_), .B(_59_), .C(_49_), .Y(_92_) );
	NAND2X1 NAND2X1_100 ( .A(A[1]), .B(B[5]), .Y(_93_) );
	INVX1 INVX1_43 ( .A(_93_), .Y(_94_) );
	AND2X2 AND2X2_15 ( .A(A[2]), .B(B[4]), .Y(_95_) );
	AND2X2 AND2X2_16 ( .A(B[3]), .B(A[3]), .Y(_96_) );
	NAND2X1 NAND2X1_101 ( .A(_95_), .B(_96_), .Y(_97_) );
	OAI21X1 OAI21X1_90 ( .A(_434_), .B(_521_), .C(_33_), .Y(_98_) );
	NAND3X1 NAND3X1_87 ( .A(_94_), .B(_98_), .C(_97_), .Y(_99_) );
	OAI21X1 OAI21X1_91 ( .A(_27_), .B(_633_), .C(_96_), .Y(_100_) );
	OAI21X1 OAI21X1_92 ( .A(_434_), .B(_521_), .C(_95_), .Y(_101_) );
	NAND3X1 NAND3X1_88 ( .A(_93_), .B(_100_), .C(_101_), .Y(_102_) );
	AND2X2 AND2X2_17 ( .A(_102_), .B(_99_), .Y(_103_) );
	AOI22X1 AOI22X1_12 ( .A(A[4]), .B(B[1]), .C(B[0]), .D(A[5]), .Y(_104_) );
	OAI21X1 OAI21X1_93 ( .A(_38_), .B(_104_), .C(_42_), .Y(_105_) );
	NAND2X1 NAND2X1_102 ( .A(A[4]), .B(B[2]), .Y(_106_) );
	INVX1 INVX1_44 ( .A(_106_), .Y(_107_) );
	AND2X2 AND2X2_18 ( .A(B[1]), .B(A[6]), .Y(_108_) );
	NAND2X1 NAND2X1_103 ( .A(_41_), .B(_108_), .Y(_109_) );
	INVX4 INVX4_5 ( .A(A[6]), .Y(_110_) );
	NAND2X1 NAND2X1_104 ( .A(B[1]), .B(A[5]), .Y(_111_) );
	OAI21X1 OAI21X1_94 ( .A(_228_), .B(_110_), .C(_111_), .Y(_112_) );
	NAND3X1 NAND3X1_89 ( .A(_107_), .B(_112_), .C(_109_), .Y(_113_) );
	NAND3X1 NAND3X1_90 ( .A(B[0]), .B(A[6]), .C(_111_), .Y(_114_) );
	NAND2X1 NAND2X1_105 ( .A(B[0]), .B(A[6]), .Y(_115_) );
	NAND3X1 NAND3X1_91 ( .A(B[1]), .B(A[5]), .C(_115_), .Y(_116_) );
	NAND3X1 NAND3X1_92 ( .A(_106_), .B(_114_), .C(_116_), .Y(_117_) );
	NAND3X1 NAND3X1_93 ( .A(_117_), .B(_105_), .C(_113_), .Y(_118_) );
	INVX1 INVX1_45 ( .A(_111_), .Y(_119_) );
	AOI22X1 AOI22X1_13 ( .A(_643_), .B(_119_), .C(_39_), .D(_44_), .Y(_120_) );
	AOI21X1 AOI21X1_61 ( .A(_114_), .B(_116_), .C(_106_), .Y(_121_) );
	AOI22X1 AOI22X1_14 ( .A(A[4]), .B(B[2]), .C(_112_), .D(_109_), .Y(_122_) );
	OAI21X1 OAI21X1_95 ( .A(_121_), .B(_122_), .C(_120_), .Y(_123_) );
	NAND3X1 NAND3X1_94 ( .A(_118_), .B(_103_), .C(_123_), .Y(_124_) );
	NAND2X1 NAND2X1_106 ( .A(_99_), .B(_102_), .Y(_125_) );
	OAI21X1 OAI21X1_96 ( .A(_121_), .B(_122_), .C(_105_), .Y(_126_) );
	NAND3X1 NAND3X1_95 ( .A(_117_), .B(_120_), .C(_113_), .Y(_127_) );
	NAND3X1 NAND3X1_96 ( .A(_125_), .B(_127_), .C(_126_), .Y(_128_) );
	NAND3X1 NAND3X1_97 ( .A(_124_), .B(_128_), .C(_92_), .Y(_129_) );
	NOR3X1 NOR3X1_7 ( .A(_50_), .B(_52_), .C(_51_), .Y(_130_) );
	AOI21X1 AOI21X1_62 ( .A(_36_), .B(_53_), .C(_130_), .Y(_131_) );
	AOI21X1 AOI21X1_63 ( .A(_126_), .B(_127_), .C(_125_), .Y(_132_) );
	AOI21X1 AOI21X1_64 ( .A(_123_), .B(_118_), .C(_103_), .Y(_133_) );
	OAI21X1 OAI21X1_97 ( .A(_132_), .B(_133_), .C(_131_), .Y(_134_) );
	NAND3X1 NAND3X1_98 ( .A(_90_), .B(_129_), .C(_134_), .Y(_135_) );
	INVX1 INVX1_46 ( .A(_90_), .Y(_136_) );
	OAI21X1 OAI21X1_98 ( .A(_132_), .B(_133_), .C(_92_), .Y(_137_) );
	NAND3X1 NAND3X1_99 ( .A(_124_), .B(_128_), .C(_131_), .Y(_138_) );
	NAND3X1 NAND3X1_100 ( .A(_136_), .B(_138_), .C(_137_), .Y(_139_) );
	NAND3X1 NAND3X1_101 ( .A(_135_), .B(_139_), .C(_84_), .Y(_140_) );
	NOR3X1 NOR3X1_8 ( .A(_66_), .B(_67_), .C(_65_), .Y(_141_) );
	AOI21X1 AOI21X1_65 ( .A(_23_), .B(_68_), .C(_141_), .Y(_142_) );
	AOI22X1 AOI22X1_15 ( .A(_87_), .B(_89_), .C(_138_), .D(_137_), .Y(_143_) );
	AOI21X1 AOI21X1_66 ( .A(_134_), .B(_129_), .C(_90_), .Y(_144_) );
	OAI21X1 OAI21X1_99 ( .A(_143_), .B(_144_), .C(_142_), .Y(_145_) );
	NAND3X1 NAND3X1_102 ( .A(_140_), .B(_82_), .C(_145_), .Y(_146_) );
	OAI21X1 OAI21X1_100 ( .A(_143_), .B(_144_), .C(_84_), .Y(_147_) );
	NAND3X1 NAND3X1_103 ( .A(_135_), .B(_139_), .C(_142_), .Y(_148_) );
	NAND3X1 NAND3X1_104 ( .A(_79_), .B(_147_), .C(_148_), .Y(_149_) );
	NAND2X1 NAND2X1_107 ( .A(_146_), .B(_149_), .Y(_150_) );
	XNOR2X1 XNOR2X1_8 ( .A(_150_), .B(_78_), .Y(_0__6_) );
	NAND3X1 NAND3X1_105 ( .A(_16_), .B(_80_), .C(_79_), .Y(_151_) );
	AOI21X1 AOI21X1_67 ( .A(_145_), .B(_140_), .C(_82_), .Y(_152_) );
	OAI21X1 OAI21X1_101 ( .A(_151_), .B(_152_), .C(_146_), .Y(_153_) );
	INVX1 INVX1_47 ( .A(_140_), .Y(_154_) );
	NAND2X1 NAND2X1_108 ( .A(_88_), .B(_86_), .Y(_155_) );
	INVX1 INVX1_48 ( .A(_155_), .Y(_156_) );
	AOI21X1 AOI21X1_68 ( .A(_124_), .B(_128_), .C(_92_), .Y(_157_) );
	OAI21X1 OAI21X1_102 ( .A(_136_), .B(_157_), .C(_129_), .Y(_158_) );
	NAND2X1 NAND2X1_109 ( .A(A[0]), .B(B[7]), .Y(_159_) );
	NOR2X1 NOR2X1_42 ( .A(_248_), .B(_85__bF_buf0), .Y(_160_) );
	NOR2X1 NOR2X1_43 ( .A(_95_), .B(_96_), .Y(_161_) );
	OAI21X1 OAI21X1_103 ( .A(_93_), .B(_161_), .C(_97_), .Y(_162_) );
	NAND2X1 NAND2X1_110 ( .A(_160_), .B(_162_), .Y(_163_) );
	AND2X2 AND2X2_19 ( .A(A[3]), .B(B[4]), .Y(_164_) );
	AOI22X1 AOI22X1_16 ( .A(_28_), .B(_164_), .C(_94_), .D(_98_), .Y(_165_) );
	OAI21X1 OAI21X1_104 ( .A(_248_), .B(_85__bF_buf3), .C(_165_), .Y(_166_) );
	NAND3X1 NAND3X1_106 ( .A(_159_), .B(_166_), .C(_163_), .Y(_167_) );
	INVX1 INVX1_49 ( .A(_159_), .Y(_168_) );
	INVX1 INVX1_50 ( .A(_160_), .Y(_169_) );
	NOR2X1 NOR2X1_44 ( .A(_169_), .B(_165_), .Y(_170_) );
	NOR2X1 NOR2X1_45 ( .A(_160_), .B(_162_), .Y(_171_) );
	OAI21X1 OAI21X1_105 ( .A(_170_), .B(_171_), .C(_168_), .Y(_172_) );
	NAND2X1 NAND2X1_111 ( .A(_167_), .B(_172_), .Y(_173_) );
	AOI21X1 AOI21X1_69 ( .A(_113_), .B(_117_), .C(_105_), .Y(_174_) );
	OAI21X1 OAI21X1_106 ( .A(_125_), .B(_174_), .C(_118_), .Y(_175_) );
	NAND2X1 NAND2X1_112 ( .A(A[2]), .B(B[5]), .Y(_176_) );
	AND2X2 AND2X2_20 ( .A(B[3]), .B(A[4]), .Y(_177_) );
	NAND2X1 NAND2X1_113 ( .A(_164_), .B(_177_), .Y(_178_) );
	OAI22X1 OAI22X1_6 ( .A(_434_), .B(_645_), .C(_521_), .D(_633_), .Y(_179_) );
	NAND3X1 NAND3X1_107 ( .A(_176_), .B(_179_), .C(_178_), .Y(_180_) );
	INVX1 INVX1_51 ( .A(_176_), .Y(_181_) );
	OAI21X1 OAI21X1_107 ( .A(_521_), .B(_633_), .C(_177_), .Y(_182_) );
	OAI21X1 OAI21X1_108 ( .A(_434_), .B(_645_), .C(_164_), .Y(_183_) );
	NAND3X1 NAND3X1_108 ( .A(_181_), .B(_182_), .C(_183_), .Y(_184_) );
	NAND2X1 NAND2X1_114 ( .A(_180_), .B(_184_), .Y(_185_) );
	AND2X2 AND2X2_21 ( .A(_111_), .B(_115_), .Y(_186_) );
	OAI21X1 OAI21X1_109 ( .A(_106_), .B(_186_), .C(_109_), .Y(_187_) );
	NAND2X1 NAND2X1_115 ( .A(B[2]), .B(A[5]), .Y(_188_) );
	INVX1 INVX1_52 ( .A(_188_), .Y(_189_) );
	AND2X2 AND2X2_22 ( .A(B[0]), .B(A[6]), .Y(_190_) );
	AND2X2 AND2X2_23 ( .A(B[1]), .B(A[7]), .Y(_191_) );
	NAND2X1 NAND2X1_116 ( .A(_190_), .B(_191_), .Y(_192_) );
	AOI22X1 AOI22X1_17 ( .A(B[0]), .B(A[7]), .C(B[1]), .D(A[6]), .Y(_193_) );
	INVX1 INVX1_53 ( .A(_193_), .Y(_194_) );
	NAND3X1 NAND3X1_109 ( .A(_189_), .B(_194_), .C(_192_), .Y(_195_) );
	NAND2X1 NAND2X1_117 ( .A(B[1]), .B(A[6]), .Y(_196_) );
	NAND3X1 NAND3X1_110 ( .A(B[0]), .B(A[7]), .C(_196_), .Y(_197_) );
	NAND2X1 NAND2X1_118 ( .A(B[0]), .B(A[7]), .Y(_198_) );
	NAND3X1 NAND3X1_111 ( .A(B[1]), .B(A[6]), .C(_198_), .Y(_199_) );
	NAND3X1 NAND3X1_112 ( .A(_188_), .B(_197_), .C(_199_), .Y(_200_) );
	NAND3X1 NAND3X1_113 ( .A(_200_), .B(_195_), .C(_187_), .Y(_201_) );
	AOI22X1 AOI22X1_18 ( .A(_41_), .B(_108_), .C(_107_), .D(_112_), .Y(_202_) );
	AOI21X1 AOI21X1_70 ( .A(_197_), .B(_199_), .C(_188_), .Y(_203_) );
	AOI22X1 AOI22X1_19 ( .A(B[2]), .B(A[5]), .C(_194_), .D(_192_), .Y(_204_) );
	OAI21X1 OAI21X1_110 ( .A(_203_), .B(_204_), .C(_202_), .Y(_205_) );
	NAND3X1 NAND3X1_114 ( .A(_185_), .B(_201_), .C(_205_), .Y(_206_) );
	NAND3X1 NAND3X1_115 ( .A(_181_), .B(_179_), .C(_178_), .Y(_207_) );
	NAND3X1 NAND3X1_116 ( .A(_176_), .B(_182_), .C(_183_), .Y(_208_) );
	NAND2X1 NAND2X1_119 ( .A(_207_), .B(_208_), .Y(_209_) );
	OAI21X1 OAI21X1_111 ( .A(_203_), .B(_204_), .C(_187_), .Y(_210_) );
	NAND3X1 NAND3X1_117 ( .A(_200_), .B(_202_), .C(_195_), .Y(_211_) );
	NAND3X1 NAND3X1_118 ( .A(_209_), .B(_211_), .C(_210_), .Y(_212_) );
	NAND3X1 NAND3X1_119 ( .A(_206_), .B(_212_), .C(_175_), .Y(_213_) );
	NOR3X1 NOR3X1_9 ( .A(_120_), .B(_121_), .C(_122_), .Y(_214_) );
	AOI21X1 AOI21X1_71 ( .A(_103_), .B(_123_), .C(_214_), .Y(_215_) );
	AOI22X1 AOI22X1_20 ( .A(_180_), .B(_184_), .C(_211_), .D(_210_), .Y(_216_) );
	AOI21X1 AOI21X1_72 ( .A(_205_), .B(_201_), .C(_185_), .Y(_217_) );
	OAI21X1 OAI21X1_112 ( .A(_216_), .B(_217_), .C(_215_), .Y(_218_) );
	NAND3X1 NAND3X1_120 ( .A(_173_), .B(_213_), .C(_218_), .Y(_219_) );
	NAND3X1 NAND3X1_121 ( .A(_168_), .B(_166_), .C(_163_), .Y(_220_) );
	OAI21X1 OAI21X1_113 ( .A(_170_), .B(_171_), .C(_159_), .Y(_221_) );
	NAND2X1 NAND2X1_120 ( .A(_220_), .B(_221_), .Y(_222_) );
	OAI21X1 OAI21X1_114 ( .A(_216_), .B(_217_), .C(_175_), .Y(_223_) );
	NAND3X1 NAND3X1_122 ( .A(_206_), .B(_212_), .C(_215_), .Y(_224_) );
	NAND3X1 NAND3X1_123 ( .A(_222_), .B(_224_), .C(_223_), .Y(_225_) );
	NAND3X1 NAND3X1_124 ( .A(_219_), .B(_158_), .C(_225_), .Y(_226_) );
	INVX1 INVX1_54 ( .A(_129_), .Y(_227_) );
	AOI21X1 AOI21X1_73 ( .A(_90_), .B(_134_), .C(_227_), .Y(_229_) );
	AOI21X1 AOI21X1_74 ( .A(_223_), .B(_224_), .C(_222_), .Y(_230_) );
	AOI21X1 AOI21X1_75 ( .A(_218_), .B(_213_), .C(_173_), .Y(_231_) );
	OAI21X1 OAI21X1_115 ( .A(_230_), .B(_231_), .C(_229_), .Y(_232_) );
	NAND3X1 NAND3X1_125 ( .A(_156_), .B(_226_), .C(_232_), .Y(_233_) );
	OAI21X1 OAI21X1_116 ( .A(_230_), .B(_231_), .C(_158_), .Y(_234_) );
	NAND3X1 NAND3X1_126 ( .A(_219_), .B(_225_), .C(_229_), .Y(_235_) );
	NAND3X1 NAND3X1_127 ( .A(_155_), .B(_234_), .C(_235_), .Y(_236_) );
	NAND3X1 NAND3X1_128 ( .A(_154_), .B(_233_), .C(_236_), .Y(_237_) );
	AOI21X1 AOI21X1_76 ( .A(_235_), .B(_234_), .C(_155_), .Y(_238_) );
	AOI21X1 AOI21X1_77 ( .A(_232_), .B(_226_), .C(_156_), .Y(_239_) );
	OAI21X1 OAI21X1_117 ( .A(_239_), .B(_238_), .C(_140_), .Y(_240_) );
	NAND2X1 NAND2X1_121 ( .A(_237_), .B(_240_), .Y(_241_) );
	XNOR2X1 XNOR2X1_9 ( .A(_241_), .B(_153_), .Y(_0__7_) );
	AOI21X1 AOI21X1_78 ( .A(_148_), .B(_147_), .C(_79_), .Y(_242_) );
	AOI21X1 AOI21X1_79 ( .A(_149_), .B(_78_), .C(_242_), .Y(_243_) );
	NOR2X1 NOR2X1_46 ( .A(_143_), .B(_144_), .Y(_244_) );
	AOI22X1 AOI22X1_21 ( .A(_84_), .B(_244_), .C(_233_), .D(_236_), .Y(_245_) );
	OAI21X1 OAI21X1_118 ( .A(_245_), .B(_243_), .C(_237_), .Y(_246_) );
	AOI21X1 AOI21X1_80 ( .A(_225_), .B(_219_), .C(_158_), .Y(_247_) );
	OAI21X1 OAI21X1_119 ( .A(_155_), .B(_247_), .C(_226_), .Y(_250_) );
	OAI21X1 OAI21X1_120 ( .A(_159_), .B(_171_), .C(_163_), .Y(_251_) );
	INVX1 INVX1_55 ( .A(_251_), .Y(_252_) );
	AOI21X1 AOI21X1_81 ( .A(_206_), .B(_212_), .C(_175_), .Y(_253_) );
	OAI21X1 OAI21X1_121 ( .A(_222_), .B(_253_), .C(_213_), .Y(_254_) );
	NAND2X1 NAND2X1_122 ( .A(A[1]), .B(B[7]), .Y(_255_) );
	NOR2X1 NOR2X1_47 ( .A(_27_), .B(_85__bF_buf2), .Y(_256_) );
	NOR2X1 NOR2X1_48 ( .A(_164_), .B(_177_), .Y(_257_) );
	OAI21X1 OAI21X1_122 ( .A(_176_), .B(_257_), .C(_178_), .Y(_258_) );
	NAND2X1 NAND2X1_123 ( .A(_256_), .B(_258_), .Y(_259_) );
	AND2X2 AND2X2_24 ( .A(A[4]), .B(B[4]), .Y(_260_) );
	AOI22X1 AOI22X1_22 ( .A(_96_), .B(_260_), .C(_181_), .D(_179_), .Y(_261_) );
	OAI21X1 OAI21X1_123 ( .A(_27_), .B(_85__bF_buf1), .C(_261_), .Y(_262_) );
	NAND3X1 NAND3X1_129 ( .A(_255_), .B(_262_), .C(_259_), .Y(_263_) );
	INVX1 INVX1_56 ( .A(_255_), .Y(_264_) );
	OAI21X1 OAI21X1_124 ( .A(_27_), .B(_85__bF_buf0), .C(_258_), .Y(_265_) );
	NAND2X1 NAND2X1_124 ( .A(_256_), .B(_261_), .Y(_266_) );
	NAND3X1 NAND3X1_130 ( .A(_264_), .B(_266_), .C(_265_), .Y(_267_) );
	AOI21X1 AOI21X1_82 ( .A(_195_), .B(_200_), .C(_187_), .Y(_268_) );
	OAI21X1 OAI21X1_125 ( .A(_209_), .B(_268_), .C(_201_), .Y(_269_) );
	NAND2X1 NAND2X1_125 ( .A(A[3]), .B(B[5]), .Y(_272_) );
	AND2X2 AND2X2_25 ( .A(B[3]), .B(A[5]), .Y(_273_) );
	NAND2X1 NAND2X1_126 ( .A(_260_), .B(_273_), .Y(_274_) );
	INVX4 INVX4_6 ( .A(A[5]), .Y(_275_) );
	NAND2X1 NAND2X1_127 ( .A(A[4]), .B(B[4]), .Y(_276_) );
	OAI21X1 OAI21X1_126 ( .A(_434_), .B(_275_), .C(_276_), .Y(_277_) );
	NAND3X1 NAND3X1_131 ( .A(_272_), .B(_277_), .C(_274_), .Y(_278_) );
	INVX1 INVX1_57 ( .A(_272_), .Y(_279_) );
endmodule
