module fir_step4 ( gnd, vdd, clk, rst, x, dataout);

input gnd, vdd;
input clk;
input rst;
input [7:0] x;
output [9:0] dataout;

	BUFX4 BUFX4_1 ( .gnd(gnd), .vdd(vdd), .A(clk), .Y(clk_bF_buf4) );
	BUFX4 BUFX4_2 ( .gnd(gnd), .vdd(vdd), .A(clk), .Y(clk_bF_buf3) );
	BUFX4 BUFX4_3 ( .gnd(gnd), .vdd(vdd), .A(clk), .Y(clk_bF_buf2) );
	BUFX4 BUFX4_4 ( .gnd(gnd), .vdd(vdd), .A(clk), .Y(clk_bF_buf1) );
	BUFX4 BUFX4_5 ( .gnd(gnd), .vdd(vdd), .A(clk), .Y(clk_bF_buf0) );
	BUFX4 BUFX4_6 ( .gnd(gnd), .vdd(vdd), .A(rst), .Y(rst_bF_buf4) );
	BUFX4 BUFX4_7 ( .gnd(gnd), .vdd(vdd), .A(rst), .Y(rst_bF_buf3) );
	BUFX4 BUFX4_8 ( .gnd(gnd), .vdd(vdd), .A(rst), .Y(rst_bF_buf2) );
	BUFX4 BUFX4_9 ( .gnd(gnd), .vdd(vdd), .A(rst), .Y(rst_bF_buf1) );
	BUFX4 BUFX4_10 ( .gnd(gnd), .vdd(vdd), .A(rst), .Y(rst_bF_buf0) );
	INVX1 INVX1_1 ( .gnd(gnd), .vdd(vdd), .A(d12_3_), .Y(_123_) );
	NAND2X1 NAND2X1_1 ( .gnd(gnd), .vdd(vdd), .A(d11_4_), .B(x[5]), .Y(_124_) );
	INVX1 INVX1_2 ( .gnd(gnd), .vdd(vdd), .A(_124_), .Y(_125_) );
	NOR2X1 NOR2X1_1 ( .gnd(gnd), .vdd(vdd), .A(d11_4_), .B(x[5]), .Y(_126_) );
	OAI21X1 OAI21X1_1 ( .gnd(gnd), .vdd(vdd), .A(_126_), .B(_125_), .C(_123_), .Y(_127_) );
	INVX1 INVX1_3 ( .gnd(gnd), .vdd(vdd), .A(_126_), .Y(_128_) );
	NAND3X1 NAND3X1_1 ( .gnd(gnd), .vdd(vdd), .A(d12_3_), .B(_124_), .C(_128_), .Y(_129_) );
	NAND3X1 NAND3X1_2 ( .gnd(gnd), .vdd(vdd), .A(d13_2_), .B(_127_), .C(_129_), .Y(_130_) );
	INVX2 INVX2_1 ( .gnd(gnd), .vdd(vdd), .A(_130_), .Y(_131_) );
	AOI21X1 AOI21X1_1 ( .gnd(gnd), .vdd(vdd), .A(_129_), .B(_127_), .C(d13_2_), .Y(_132_) );
	NOR2X1 NOR2X1_2 ( .gnd(gnd), .vdd(vdd), .A(_132_), .B(_131_), .Y(_133_) );
	NAND2X1 NAND2X1_2 ( .gnd(gnd), .vdd(vdd), .A(d14_1_), .B(_133_), .Y(_134_) );
	INVX1 INVX1_4 ( .gnd(gnd), .vdd(vdd), .A(_134_), .Y(_135_) );
	NOR2X1 NOR2X1_3 ( .gnd(gnd), .vdd(vdd), .A(d14_1_), .B(_133_), .Y(_136_) );
	NOR2X1 NOR2X1_4 ( .gnd(gnd), .vdd(vdd), .A(_136_), .B(_135_), .Y(_187__0_) );
	OAI21X1 OAI21X1_2 ( .gnd(gnd), .vdd(vdd), .A(_123_), .B(_126_), .C(_124_), .Y(_137_) );
	INVX1 INVX1_5 ( .gnd(gnd), .vdd(vdd), .A(d12_4_), .Y(_138_) );
	AND2X2 AND2X2_1 ( .gnd(gnd), .vdd(vdd), .A(d11_5_), .B(x[6]), .Y(_139_) );
	NOR2X1 NOR2X1_5 ( .gnd(gnd), .vdd(vdd), .A(d11_5_), .B(x[6]), .Y(_140_) );
	OAI21X1 OAI21X1_3 ( .gnd(gnd), .vdd(vdd), .A(_140_), .B(_139_), .C(_138_), .Y(_141_) );
	NAND2X1 NAND2X1_3 ( .gnd(gnd), .vdd(vdd), .A(d11_5_), .B(x[6]), .Y(_142_) );
	OR2X2 OR2X2_1 ( .gnd(gnd), .vdd(vdd), .A(d11_5_), .B(x[6]), .Y(_143_) );
	NAND3X1 NAND3X1_3 ( .gnd(gnd), .vdd(vdd), .A(d12_4_), .B(_142_), .C(_143_), .Y(_144_) );
	NAND3X1 NAND3X1_4 ( .gnd(gnd), .vdd(vdd), .A(_137_), .B(_141_), .C(_144_), .Y(_145_) );
	INVX1 INVX1_6 ( .gnd(gnd), .vdd(vdd), .A(_137_), .Y(_146_) );
	NAND2X1 NAND2X1_4 ( .gnd(gnd), .vdd(vdd), .A(_141_), .B(_144_), .Y(_147_) );
	NAND2X1 NAND2X1_5 ( .gnd(gnd), .vdd(vdd), .A(_146_), .B(_147_), .Y(_148_) );
	NAND3X1 NAND3X1_5 ( .gnd(gnd), .vdd(vdd), .A(d13_3_), .B(_145_), .C(_148_), .Y(_149_) );
	INVX1 INVX1_7 ( .gnd(gnd), .vdd(vdd), .A(d13_3_), .Y(_150_) );
	NAND2X1 NAND2X1_6 ( .gnd(gnd), .vdd(vdd), .A(_137_), .B(_147_), .Y(_151_) );
	NAND3X1 NAND3X1_6 ( .gnd(gnd), .vdd(vdd), .A(_141_), .B(_144_), .C(_146_), .Y(_152_) );
	NAND3X1 NAND3X1_7 ( .gnd(gnd), .vdd(vdd), .A(_150_), .B(_152_), .C(_151_), .Y(_153_) );
	NAND3X1 NAND3X1_8 ( .gnd(gnd), .vdd(vdd), .A(_130_), .B(_149_), .C(_153_), .Y(_154_) );
	INVX1 INVX1_8 ( .gnd(gnd), .vdd(vdd), .A(_145_), .Y(_155_) );
	AOI21X1 AOI21X1_2 ( .gnd(gnd), .vdd(vdd), .A(_144_), .B(_141_), .C(_137_), .Y(_156_) );
	OAI21X1 OAI21X1_4 ( .gnd(gnd), .vdd(vdd), .A(_156_), .B(_155_), .C(d13_3_), .Y(_157_) );
	NAND3X1 NAND3X1_9 ( .gnd(gnd), .vdd(vdd), .A(_150_), .B(_145_), .C(_148_), .Y(_158_) );
	NAND3X1 NAND3X1_10 ( .gnd(gnd), .vdd(vdd), .A(_131_), .B(_158_), .C(_157_), .Y(_159_) );
	NAND3X1 NAND3X1_11 ( .gnd(gnd), .vdd(vdd), .A(d14_2_), .B(_154_), .C(_159_), .Y(_160_) );
	INVX1 INVX1_9 ( .gnd(gnd), .vdd(vdd), .A(d14_2_), .Y(_161_) );
	NAND3X1 NAND3X1_12 ( .gnd(gnd), .vdd(vdd), .A(_131_), .B(_149_), .C(_153_), .Y(_162_) );
	NAND3X1 NAND3X1_13 ( .gnd(gnd), .vdd(vdd), .A(_130_), .B(_158_), .C(_157_), .Y(_163_) );
	NAND3X1 NAND3X1_14 ( .gnd(gnd), .vdd(vdd), .A(_161_), .B(_162_), .C(_163_), .Y(_164_) );
	AOI21X1 AOI21X1_3 ( .gnd(gnd), .vdd(vdd), .A(_160_), .B(_164_), .C(_134_), .Y(_165_) );
	NAND2X1 NAND2X1_7 ( .gnd(gnd), .vdd(vdd), .A(_160_), .B(_164_), .Y(_166_) );
	NOR2X1 NOR2X1_6 ( .gnd(gnd), .vdd(vdd), .A(_135_), .B(_166_), .Y(_167_) );
	NOR2X1 NOR2X1_7 ( .gnd(gnd), .vdd(vdd), .A(_165_), .B(_167_), .Y(_187__1_) );
	AOI21X1 AOI21X1_4 ( .gnd(gnd), .vdd(vdd), .A(_149_), .B(_153_), .C(_131_), .Y(_168_) );
	OAI21X1 OAI21X1_5 ( .gnd(gnd), .vdd(vdd), .A(_161_), .B(_168_), .C(_162_), .Y(_169_) );
	OAI21X1 OAI21X1_6 ( .gnd(gnd), .vdd(vdd), .A(_150_), .B(_156_), .C(_145_), .Y(_170_) );
	INVX1 INVX1_10 ( .gnd(gnd), .vdd(vdd), .A(d13_4_), .Y(_171_) );
	OAI21X1 OAI21X1_7 ( .gnd(gnd), .vdd(vdd), .A(_138_), .B(_140_), .C(_142_), .Y(_172_) );
	NAND2X1 NAND2X1_8 ( .gnd(gnd), .vdd(vdd), .A(d11_6_), .B(x[7]), .Y(_173_) );
	OR2X2 OR2X2_2 ( .gnd(gnd), .vdd(vdd), .A(d11_6_), .B(x[7]), .Y(_174_) );
	AOI21X1 AOI21X1_5 ( .gnd(gnd), .vdd(vdd), .A(_174_), .B(_173_), .C(d12_5_), .Y(_175_) );
	INVX1 INVX1_11 ( .gnd(gnd), .vdd(vdd), .A(d12_5_), .Y(_176_) );
	AND2X2 AND2X2_2 ( .gnd(gnd), .vdd(vdd), .A(d11_6_), .B(x[7]), .Y(_177_) );
	NOR2X1 NOR2X1_8 ( .gnd(gnd), .vdd(vdd), .A(d11_6_), .B(x[7]), .Y(_178_) );
	NOR3X1 NOR3X1_1 ( .gnd(gnd), .vdd(vdd), .A(_176_), .B(_178_), .C(_177_), .Y(_179_) );
	OAI21X1 OAI21X1_8 ( .gnd(gnd), .vdd(vdd), .A(_175_), .B(_179_), .C(_172_), .Y(_180_) );
	AOI21X1 AOI21X1_6 ( .gnd(gnd), .vdd(vdd), .A(_143_), .B(d12_4_), .C(_139_), .Y(_181_) );
	OAI21X1 OAI21X1_9 ( .gnd(gnd), .vdd(vdd), .A(_178_), .B(_177_), .C(_176_), .Y(_182_) );
	NAND3X1 NAND3X1_15 ( .gnd(gnd), .vdd(vdd), .A(d12_5_), .B(_173_), .C(_174_), .Y(_183_) );
	NAND3X1 NAND3X1_16 ( .gnd(gnd), .vdd(vdd), .A(_182_), .B(_183_), .C(_181_), .Y(_184_) );
	NAND3X1 NAND3X1_17 ( .gnd(gnd), .vdd(vdd), .A(_171_), .B(_184_), .C(_180_), .Y(_185_) );
	NAND3X1 NAND3X1_18 ( .gnd(gnd), .vdd(vdd), .A(_172_), .B(_182_), .C(_183_), .Y(_186_) );
	OAI21X1 OAI21X1_10 ( .gnd(gnd), .vdd(vdd), .A(_175_), .B(_179_), .C(_181_), .Y(_0_) );
	NAND3X1 NAND3X1_19 ( .gnd(gnd), .vdd(vdd), .A(d13_4_), .B(_186_), .C(_0_), .Y(_1_) );
	NAND3X1 NAND3X1_20 ( .gnd(gnd), .vdd(vdd), .A(_170_), .B(_185_), .C(_1_), .Y(_2_) );
	AOI21X1 AOI21X1_7 ( .gnd(gnd), .vdd(vdd), .A(_148_), .B(d13_3_), .C(_155_), .Y(_3_) );
	AOI21X1 AOI21X1_8 ( .gnd(gnd), .vdd(vdd), .A(_0_), .B(_186_), .C(d13_4_), .Y(_4_) );
	AOI21X1 AOI21X1_9 ( .gnd(gnd), .vdd(vdd), .A(_180_), .B(_184_), .C(_171_), .Y(_5_) );
	OAI21X1 OAI21X1_11 ( .gnd(gnd), .vdd(vdd), .A(_4_), .B(_5_), .C(_3_), .Y(_6_) );
	AOI21X1 AOI21X1_10 ( .gnd(gnd), .vdd(vdd), .A(_6_), .B(_2_), .C(d14_3_), .Y(_7_) );
	INVX1 INVX1_12 ( .gnd(gnd), .vdd(vdd), .A(d14_3_), .Y(_8_) );
	OAI21X1 OAI21X1_12 ( .gnd(gnd), .vdd(vdd), .A(_4_), .B(_5_), .C(_170_), .Y(_9_) );
	NAND3X1 NAND3X1_21 ( .gnd(gnd), .vdd(vdd), .A(_185_), .B(_1_), .C(_3_), .Y(_10_) );
	AOI21X1 AOI21X1_11 ( .gnd(gnd), .vdd(vdd), .A(_9_), .B(_10_), .C(_8_), .Y(_11_) );
	OAI21X1 OAI21X1_13 ( .gnd(gnd), .vdd(vdd), .A(_7_), .B(_11_), .C(_169_), .Y(_12_) );
	AOI21X1 AOI21X1_12 ( .gnd(gnd), .vdd(vdd), .A(_157_), .B(_158_), .C(_130_), .Y(_13_) );
	AOI21X1 AOI21X1_13 ( .gnd(gnd), .vdd(vdd), .A(d14_2_), .B(_163_), .C(_13_), .Y(_14_) );
	NAND3X1 NAND3X1_22 ( .gnd(gnd), .vdd(vdd), .A(_8_), .B(_10_), .C(_9_), .Y(_15_) );
	NAND3X1 NAND3X1_23 ( .gnd(gnd), .vdd(vdd), .A(d14_3_), .B(_2_), .C(_6_), .Y(_16_) );
	NAND3X1 NAND3X1_24 ( .gnd(gnd), .vdd(vdd), .A(_16_), .B(_15_), .C(_14_), .Y(_17_) );
	NAND2X1 NAND2X1_9 ( .gnd(gnd), .vdd(vdd), .A(_17_), .B(_12_), .Y(_18_) );
	XOR2X1 XOR2X1_1 ( .gnd(gnd), .vdd(vdd), .A(_18_), .B(_165_), .Y(_187__2_) );
	NAND3X1 NAND3X1_25 ( .gnd(gnd), .vdd(vdd), .A(_16_), .B(_15_), .C(_169_), .Y(_19_) );
	OAI21X1 OAI21X1_14 ( .gnd(gnd), .vdd(vdd), .A(_7_), .B(_11_), .C(_14_), .Y(_20_) );
	NAND3X1 NAND3X1_26 ( .gnd(gnd), .vdd(vdd), .A(_165_), .B(_19_), .C(_20_), .Y(_21_) );
	NAND2X1 NAND2X1_10 ( .gnd(gnd), .vdd(vdd), .A(_19_), .B(_21_), .Y(_22_) );
	AOI21X1 AOI21X1_14 ( .gnd(gnd), .vdd(vdd), .A(_185_), .B(_1_), .C(_170_), .Y(_23_) );
	OAI21X1 OAI21X1_15 ( .gnd(gnd), .vdd(vdd), .A(_8_), .B(_23_), .C(_2_), .Y(_24_) );
	AOI21X1 AOI21X1_15 ( .gnd(gnd), .vdd(vdd), .A(_183_), .B(_182_), .C(_172_), .Y(_25_) );
	OAI21X1 OAI21X1_16 ( .gnd(gnd), .vdd(vdd), .A(_171_), .B(_25_), .C(_186_), .Y(_26_) );
	INVX1 INVX1_13 ( .gnd(gnd), .vdd(vdd), .A(d14_4_), .Y(_27_) );
	OAI21X1 OAI21X1_17 ( .gnd(gnd), .vdd(vdd), .A(_176_), .B(_178_), .C(_173_), .Y(_28_) );
	INVX1 INVX1_14 ( .gnd(gnd), .vdd(vdd), .A(d13_5_), .Y(_29_) );
	NOR2X1 NOR2X1_9 ( .gnd(gnd), .vdd(vdd), .A(d12_6_), .B(d11_7_), .Y(_30_) );
	AND2X2 AND2X2_3 ( .gnd(gnd), .vdd(vdd), .A(d12_6_), .B(d11_7_), .Y(_31_) );
	NOR3X1 NOR3X1_2 ( .gnd(gnd), .vdd(vdd), .A(_29_), .B(_30_), .C(_31_), .Y(_32_) );
	OR2X2 OR2X2_3 ( .gnd(gnd), .vdd(vdd), .A(d12_6_), .B(d11_7_), .Y(_33_) );
	NAND2X1 NAND2X1_11 ( .gnd(gnd), .vdd(vdd), .A(d12_6_), .B(d11_7_), .Y(_34_) );
	AOI21X1 AOI21X1_16 ( .gnd(gnd), .vdd(vdd), .A(_33_), .B(_34_), .C(d13_5_), .Y(_35_) );
	OAI21X1 OAI21X1_18 ( .gnd(gnd), .vdd(vdd), .A(_35_), .B(_32_), .C(_28_), .Y(_36_) );
	INVX1 INVX1_15 ( .gnd(gnd), .vdd(vdd), .A(_28_), .Y(_37_) );
	NAND3X1 NAND3X1_27 ( .gnd(gnd), .vdd(vdd), .A(d13_5_), .B(_34_), .C(_33_), .Y(_38_) );
	OAI21X1 OAI21X1_19 ( .gnd(gnd), .vdd(vdd), .A(_30_), .B(_31_), .C(_29_), .Y(_39_) );
	NAND3X1 NAND3X1_28 ( .gnd(gnd), .vdd(vdd), .A(_38_), .B(_39_), .C(_37_), .Y(_40_) );
	NAND3X1 NAND3X1_29 ( .gnd(gnd), .vdd(vdd), .A(_27_), .B(_36_), .C(_40_), .Y(_41_) );
	NAND3X1 NAND3X1_30 ( .gnd(gnd), .vdd(vdd), .A(_28_), .B(_39_), .C(_38_), .Y(_42_) );
	OAI21X1 OAI21X1_20 ( .gnd(gnd), .vdd(vdd), .A(_35_), .B(_32_), .C(_37_), .Y(_43_) );
	NAND3X1 NAND3X1_31 ( .gnd(gnd), .vdd(vdd), .A(d14_4_), .B(_42_), .C(_43_), .Y(_44_) );
	NAND3X1 NAND3X1_32 ( .gnd(gnd), .vdd(vdd), .A(_26_), .B(_44_), .C(_41_), .Y(_45_) );
	INVX1 INVX1_16 ( .gnd(gnd), .vdd(vdd), .A(_186_), .Y(_46_) );
	AOI21X1 AOI21X1_17 ( .gnd(gnd), .vdd(vdd), .A(d13_4_), .B(_0_), .C(_46_), .Y(_47_) );
	AOI21X1 AOI21X1_18 ( .gnd(gnd), .vdd(vdd), .A(_43_), .B(_42_), .C(d14_4_), .Y(_48_) );
	AOI21X1 AOI21X1_19 ( .gnd(gnd), .vdd(vdd), .A(_40_), .B(_36_), .C(_27_), .Y(_49_) );
	OAI21X1 OAI21X1_21 ( .gnd(gnd), .vdd(vdd), .A(_48_), .B(_49_), .C(_47_), .Y(_50_) );
	NAND2X1 NAND2X1_12 ( .gnd(gnd), .vdd(vdd), .A(_45_), .B(_50_), .Y(_51_) );
	XOR2X1 XOR2X1_2 ( .gnd(gnd), .vdd(vdd), .A(_24_), .B(_51_), .Y(_52_) );
	XNOR2X1 XNOR2X1_1 ( .gnd(gnd), .vdd(vdd), .A(_22_), .B(_52_), .Y(_187__3_) );
	XNOR2X1 XNOR2X1_2 ( .gnd(gnd), .vdd(vdd), .A(_24_), .B(_51_), .Y(_53_) );
	NAND3X1 NAND3X1_33 ( .gnd(gnd), .vdd(vdd), .A(_165_), .B(_53_), .C(_18_), .Y(_54_) );
	NAND3X1 NAND3X1_34 ( .gnd(gnd), .vdd(vdd), .A(_45_), .B(_50_), .C(_24_), .Y(_55_) );
	AOI21X1 AOI21X1_20 ( .gnd(gnd), .vdd(vdd), .A(_45_), .B(_50_), .C(_24_), .Y(_56_) );
	OAI21X1 OAI21X1_22 ( .gnd(gnd), .vdd(vdd), .A(_56_), .B(_19_), .C(_55_), .Y(_57_) );
	INVX1 INVX1_17 ( .gnd(gnd), .vdd(vdd), .A(_57_), .Y(_58_) );
	NAND2X1 NAND2X1_13 ( .gnd(gnd), .vdd(vdd), .A(_42_), .B(_44_), .Y(_59_) );
	OAI21X1 OAI21X1_23 ( .gnd(gnd), .vdd(vdd), .A(_29_), .B(_30_), .C(_34_), .Y(_60_) );
	INVX1 INVX1_18 ( .gnd(gnd), .vdd(vdd), .A(d14_5_), .Y(_61_) );
	NOR2X1 NOR2X1_10 ( .gnd(gnd), .vdd(vdd), .A(d13_6_), .B(d12_7_), .Y(_62_) );
	NAND2X1 NAND2X1_14 ( .gnd(gnd), .vdd(vdd), .A(d13_6_), .B(d12_7_), .Y(_63_) );
	INVX1 INVX1_19 ( .gnd(gnd), .vdd(vdd), .A(_63_), .Y(_64_) );
	NOR2X1 NOR2X1_11 ( .gnd(gnd), .vdd(vdd), .A(_62_), .B(_64_), .Y(_65_) );
	XNOR2X1 XNOR2X1_3 ( .gnd(gnd), .vdd(vdd), .A(_65_), .B(_61_), .Y(_66_) );
	XOR2X1 XOR2X1_3 ( .gnd(gnd), .vdd(vdd), .A(_66_), .B(_60_), .Y(_67_) );
	AND2X2 AND2X2_4 ( .gnd(gnd), .vdd(vdd), .A(_67_), .B(_59_), .Y(_68_) );
	NOR2X1 NOR2X1_12 ( .gnd(gnd), .vdd(vdd), .A(_59_), .B(_67_), .Y(_69_) );
	OAI21X1 OAI21X1_24 ( .gnd(gnd), .vdd(vdd), .A(_69_), .B(_68_), .C(_45_), .Y(_70_) );
	NOR3X1 NOR3X1_3 ( .gnd(gnd), .vdd(vdd), .A(_45_), .B(_69_), .C(_68_), .Y(_71_) );
	INVX2 INVX2_2 ( .gnd(gnd), .vdd(vdd), .A(_71_), .Y(_72_) );
	NAND2X1 NAND2X1_15 ( .gnd(gnd), .vdd(vdd), .A(_70_), .B(_72_), .Y(_73_) );
	AOI21X1 AOI21X1_21 ( .gnd(gnd), .vdd(vdd), .A(_54_), .B(_58_), .C(_73_), .Y(_74_) );
	OAI21X1 OAI21X1_25 ( .gnd(gnd), .vdd(vdd), .A(_21_), .B(_52_), .C(_58_), .Y(_75_) );
	INVX1 INVX1_20 ( .gnd(gnd), .vdd(vdd), .A(_45_), .Y(_76_) );
	NAND2X1 NAND2X1_16 ( .gnd(gnd), .vdd(vdd), .A(_59_), .B(_67_), .Y(_77_) );
	INVX1 INVX1_21 ( .gnd(gnd), .vdd(vdd), .A(_69_), .Y(_78_) );
	AOI21X1 AOI21X1_22 ( .gnd(gnd), .vdd(vdd), .A(_78_), .B(_77_), .C(_76_), .Y(_79_) );
	NOR2X1 NOR2X1_13 ( .gnd(gnd), .vdd(vdd), .A(_71_), .B(_79_), .Y(_80_) );
	NOR2X1 NOR2X1_14 ( .gnd(gnd), .vdd(vdd), .A(_80_), .B(_75_), .Y(_81_) );
	NOR2X1 NOR2X1_15 ( .gnd(gnd), .vdd(vdd), .A(_74_), .B(_81_), .Y(_187__4_) );
	OAI21X1 OAI21X1_26 ( .gnd(gnd), .vdd(vdd), .A(_31_), .B(_32_), .C(_66_), .Y(_82_) );
	OAI21X1 OAI21X1_27 ( .gnd(gnd), .vdd(vdd), .A(_61_), .B(_62_), .C(_63_), .Y(_83_) );
	NAND2X1 NAND2X1_17 ( .gnd(gnd), .vdd(vdd), .A(d14_6_), .B(d13_7_), .Y(_84_) );
	INVX1 INVX1_22 ( .gnd(gnd), .vdd(vdd), .A(d14_6_), .Y(_85_) );
	INVX1 INVX1_23 ( .gnd(gnd), .vdd(vdd), .A(d13_7_), .Y(_86_) );
	NAND2X1 NAND2X1_18 ( .gnd(gnd), .vdd(vdd), .A(_85_), .B(_86_), .Y(_87_) );
	NAND2X1 NAND2X1_19 ( .gnd(gnd), .vdd(vdd), .A(_84_), .B(_87_), .Y(_88_) );
	XNOR2X1 XNOR2X1_4 ( .gnd(gnd), .vdd(vdd), .A(_88_), .B(_83_), .Y(_89_) );
	INVX1 INVX1_24 ( .gnd(gnd), .vdd(vdd), .A(_89_), .Y(_90_) );
	NAND2X1 NAND2X1_20 ( .gnd(gnd), .vdd(vdd), .A(_90_), .B(_82_), .Y(_91_) );
	NAND3X1 NAND3X1_35 ( .gnd(gnd), .vdd(vdd), .A(_60_), .B(_66_), .C(_89_), .Y(_92_) );
	NAND2X1 NAND2X1_21 ( .gnd(gnd), .vdd(vdd), .A(_92_), .B(_91_), .Y(_93_) );
	NAND2X1 NAND2X1_22 ( .gnd(gnd), .vdd(vdd), .A(_93_), .B(_77_), .Y(_94_) );
	INVX1 INVX1_25 ( .gnd(gnd), .vdd(vdd), .A(_93_), .Y(_95_) );
	NAND2X1 NAND2X1_23 ( .gnd(gnd), .vdd(vdd), .A(_68_), .B(_95_), .Y(_96_) );
	NAND2X1 NAND2X1_24 ( .gnd(gnd), .vdd(vdd), .A(_94_), .B(_96_), .Y(_97_) );
	OAI21X1 OAI21X1_28 ( .gnd(gnd), .vdd(vdd), .A(_71_), .B(_74_), .C(_97_), .Y(_98_) );
	NOR2X1 NOR2X1_16 ( .gnd(gnd), .vdd(vdd), .A(_52_), .B(_21_), .Y(_99_) );
	OAI21X1 OAI21X1_29 ( .gnd(gnd), .vdd(vdd), .A(_57_), .B(_99_), .C(_80_), .Y(_100_) );
	AND2X2 AND2X2_5 ( .gnd(gnd), .vdd(vdd), .A(_96_), .B(_94_), .Y(_101_) );
	NAND3X1 NAND3X1_36 ( .gnd(gnd), .vdd(vdd), .A(_72_), .B(_101_), .C(_100_), .Y(_102_) );
	NAND2X1 NAND2X1_25 ( .gnd(gnd), .vdd(vdd), .A(_102_), .B(_98_), .Y(_187__5_) );
	NOR3X1 NOR3X1_4 ( .gnd(gnd), .vdd(vdd), .A(_71_), .B(_79_), .C(_97_), .Y(_103_) );
	OAI21X1 OAI21X1_30 ( .gnd(gnd), .vdd(vdd), .A(_57_), .B(_99_), .C(_103_), .Y(_104_) );
	OAI21X1 OAI21X1_31 ( .gnd(gnd), .vdd(vdd), .A(_97_), .B(_72_), .C(_96_), .Y(_105_) );
	INVX1 INVX1_26 ( .gnd(gnd), .vdd(vdd), .A(_105_), .Y(_106_) );
	INVX1 INVX1_27 ( .gnd(gnd), .vdd(vdd), .A(d14_7_), .Y(_107_) );
	OAI21X1 OAI21X1_32 ( .gnd(gnd), .vdd(vdd), .A(_85_), .B(_86_), .C(_107_), .Y(_108_) );
	OR2X2 OR2X2_4 ( .gnd(gnd), .vdd(vdd), .A(_84_), .B(_107_), .Y(_109_) );
	NAND2X1 NAND2X1_26 ( .gnd(gnd), .vdd(vdd), .A(_108_), .B(_109_), .Y(_110_) );
	NAND3X1 NAND3X1_37 ( .gnd(gnd), .vdd(vdd), .A(_84_), .B(_87_), .C(_83_), .Y(_111_) );
	OAI21X1 OAI21X1_33 ( .gnd(gnd), .vdd(vdd), .A(_90_), .B(_82_), .C(_111_), .Y(_112_) );
	XNOR2X1 XNOR2X1_5 ( .gnd(gnd), .vdd(vdd), .A(_112_), .B(_110_), .Y(_113_) );
	NAND3X1 NAND3X1_38 ( .gnd(gnd), .vdd(vdd), .A(_106_), .B(_113_), .C(_104_), .Y(_114_) );
	NAND3X1 NAND3X1_39 ( .gnd(gnd), .vdd(vdd), .A(_70_), .B(_72_), .C(_101_), .Y(_115_) );
	AOI21X1 AOI21X1_23 ( .gnd(gnd), .vdd(vdd), .A(_54_), .B(_58_), .C(_115_), .Y(_116_) );
	INVX1 INVX1_28 ( .gnd(gnd), .vdd(vdd), .A(_113_), .Y(_117_) );
	OAI21X1 OAI21X1_34 ( .gnd(gnd), .vdd(vdd), .A(_105_), .B(_116_), .C(_117_), .Y(_118_) );
	NAND2X1 NAND2X1_27 ( .gnd(gnd), .vdd(vdd), .A(_114_), .B(_118_), .Y(_187__6_) );
	OAI21X1 OAI21X1_35 ( .gnd(gnd), .vdd(vdd), .A(_105_), .B(_116_), .C(_113_), .Y(_119_) );
	OAI21X1 OAI21X1_36 ( .gnd(gnd), .vdd(vdd), .A(_110_), .B(_111_), .C(_109_), .Y(_120_) );
	NOR2X1 NOR2X1_17 ( .gnd(gnd), .vdd(vdd), .A(_110_), .B(_92_), .Y(_121_) );
	NOR2X1 NOR2X1_18 ( .gnd(gnd), .vdd(vdd), .A(_120_), .B(_121_), .Y(_122_) );
	NAND2X1 NAND2X1_28 ( .gnd(gnd), .vdd(vdd), .A(_122_), .B(_119_), .Y(_187__7_) );
	BUFX2 BUFX2_1 ( .gnd(gnd), .vdd(vdd), .A(_187__0_), .Y(dataout[0]) );
	BUFX2 BUFX2_2 ( .gnd(gnd), .vdd(vdd), .A(_187__1_), .Y(dataout[1]) );
	BUFX2 BUFX2_3 ( .gnd(gnd), .vdd(vdd), .A(_187__2_), .Y(dataout[2]) );
	BUFX2 BUFX2_4 ( .gnd(gnd), .vdd(vdd), .A(_187__3_), .Y(dataout[3]) );
	BUFX2 BUFX2_5 ( .gnd(gnd), .vdd(vdd), .A(_187__4_), .Y(dataout[4]) );
	BUFX2 BUFX2_6 ( .gnd(gnd), .vdd(vdd), .A(_187__5_), .Y(dataout[5]) );
	BUFX2 BUFX2_7 ( .gnd(gnd), .vdd(vdd), .A(_187__6_), .Y(dataout[6]) );
	BUFX2 BUFX2_8 ( .gnd(gnd), .vdd(vdd), .A(_187__7_), .Y(dataout[7]) );
	BUFX2 BUFX2_9 ( .gnd(gnd), .vdd(vdd), .A(gnd), .Y(dataout[8]) );
	BUFX2 BUFX2_10 ( .gnd(gnd), .vdd(vdd), .A(gnd), .Y(dataout[9]) );
	INVX1 INVX1_29 ( .gnd(gnd), .vdd(vdd), .A(x[1]), .Y(_189_) );
	NOR2X1 NOR2X1_19 ( .gnd(gnd), .vdd(vdd), .A(rst_bF_buf4), .B(_189_), .Y(_188__1_) );
	INVX1 INVX1_30 ( .gnd(gnd), .vdd(vdd), .A(x[2]), .Y(_190_) );
	NOR2X1 NOR2X1_20 ( .gnd(gnd), .vdd(vdd), .A(rst_bF_buf3), .B(_190_), .Y(_188__2_) );
	INVX1 INVX1_31 ( .gnd(gnd), .vdd(vdd), .A(x[3]), .Y(_191_) );
	NOR2X1 NOR2X1_21 ( .gnd(gnd), .vdd(vdd), .A(rst_bF_buf2), .B(_191_), .Y(_188__3_) );
	INVX1 INVX1_32 ( .gnd(gnd), .vdd(vdd), .A(x[4]), .Y(_192_) );
	NOR2X1 NOR2X1_22 ( .gnd(gnd), .vdd(vdd), .A(rst_bF_buf1), .B(_192_), .Y(_188__4_) );
	INVX1 INVX1_33 ( .gnd(gnd), .vdd(vdd), .A(x[5]), .Y(_193_) );
	NOR2X1 NOR2X1_23 ( .gnd(gnd), .vdd(vdd), .A(rst_bF_buf0), .B(_193_), .Y(_188__5_) );
	INVX1 INVX1_34 ( .gnd(gnd), .vdd(vdd), .A(x[6]), .Y(_194_) );
	NOR2X1 NOR2X1_24 ( .gnd(gnd), .vdd(vdd), .A(rst_bF_buf4), .B(_194_), .Y(_188__6_) );
	INVX1 INVX1_35 ( .gnd(gnd), .vdd(vdd), .A(x[7]), .Y(_195_) );
	NOR2X1 NOR2X1_25 ( .gnd(gnd), .vdd(vdd), .A(rst_bF_buf3), .B(_195_), .Y(_188__7_) );
	DFFPOSX1 DFFPOSX1_1 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf4), .D(_188__1_), .Q(d11_1_) );
	DFFPOSX1 DFFPOSX1_2 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf3), .D(_188__2_), .Q(d11_2_) );
	DFFPOSX1 DFFPOSX1_3 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf2), .D(_188__3_), .Q(d11_3_) );
	DFFPOSX1 DFFPOSX1_4 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf1), .D(_188__4_), .Q(d11_4_) );
	DFFPOSX1 DFFPOSX1_5 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf0), .D(_188__5_), .Q(d11_5_) );
	DFFPOSX1 DFFPOSX1_6 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf4), .D(_188__6_), .Q(d11_6_) );
	DFFPOSX1 DFFPOSX1_7 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf3), .D(_188__7_), .Q(d11_7_) );
	INVX1 INVX1_36 ( .gnd(gnd), .vdd(vdd), .A(d11_1_), .Y(_197_) );
	NOR2X1 NOR2X1_26 ( .gnd(gnd), .vdd(vdd), .A(rst_bF_buf2), .B(_197_), .Y(_196__1_) );
	INVX1 INVX1_37 ( .gnd(gnd), .vdd(vdd), .A(d11_2_), .Y(_198_) );
	NOR2X1 NOR2X1_27 ( .gnd(gnd), .vdd(vdd), .A(rst_bF_buf1), .B(_198_), .Y(_196__2_) );
	INVX1 INVX1_38 ( .gnd(gnd), .vdd(vdd), .A(d11_3_), .Y(_199_) );
	NOR2X1 NOR2X1_28 ( .gnd(gnd), .vdd(vdd), .A(rst_bF_buf0), .B(_199_), .Y(_196__3_) );
	INVX1 INVX1_39 ( .gnd(gnd), .vdd(vdd), .A(d11_4_), .Y(_200_) );
	NOR2X1 NOR2X1_29 ( .gnd(gnd), .vdd(vdd), .A(rst_bF_buf4), .B(_200_), .Y(_196__4_) );
	INVX1 INVX1_40 ( .gnd(gnd), .vdd(vdd), .A(d11_5_), .Y(_201_) );
	NOR2X1 NOR2X1_30 ( .gnd(gnd), .vdd(vdd), .A(rst_bF_buf3), .B(_201_), .Y(_196__5_) );
	INVX1 INVX1_41 ( .gnd(gnd), .vdd(vdd), .A(d11_6_), .Y(_202_) );
	NOR2X1 NOR2X1_31 ( .gnd(gnd), .vdd(vdd), .A(rst_bF_buf2), .B(_202_), .Y(_196__6_) );
	INVX1 INVX1_42 ( .gnd(gnd), .vdd(vdd), .A(d11_7_), .Y(_203_) );
	NOR2X1 NOR2X1_32 ( .gnd(gnd), .vdd(vdd), .A(rst_bF_buf1), .B(_203_), .Y(_196__7_) );
	DFFPOSX1 DFFPOSX1_8 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf2), .D(_196__1_), .Q(d12_1_) );
	DFFPOSX1 DFFPOSX1_9 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf1), .D(_196__2_), .Q(d12_2_) );
	DFFPOSX1 DFFPOSX1_10 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf0), .D(_196__3_), .Q(d12_3_) );
	DFFPOSX1 DFFPOSX1_11 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf4), .D(_196__4_), .Q(d12_4_) );
	DFFPOSX1 DFFPOSX1_12 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf3), .D(_196__5_), .Q(d12_5_) );
	DFFPOSX1 DFFPOSX1_13 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf2), .D(_196__6_), .Q(d12_6_) );
	DFFPOSX1 DFFPOSX1_14 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf1), .D(_196__7_), .Q(d12_7_) );
	INVX1 INVX1_43 ( .gnd(gnd), .vdd(vdd), .A(d12_1_), .Y(_205_) );
	NOR2X1 NOR2X1_33 ( .gnd(gnd), .vdd(vdd), .A(rst_bF_buf0), .B(_205_), .Y(_204__1_) );
	INVX1 INVX1_44 ( .gnd(gnd), .vdd(vdd), .A(d12_2_), .Y(_206_) );
	NOR2X1 NOR2X1_34 ( .gnd(gnd), .vdd(vdd), .A(rst_bF_buf4), .B(_206_), .Y(_204__2_) );
	INVX1 INVX1_45 ( .gnd(gnd), .vdd(vdd), .A(d12_3_), .Y(_207_) );
	NOR2X1 NOR2X1_35 ( .gnd(gnd), .vdd(vdd), .A(rst_bF_buf3), .B(_207_), .Y(_204__3_) );
	INVX1 INVX1_46 ( .gnd(gnd), .vdd(vdd), .A(d12_4_), .Y(_208_) );
	NOR2X1 NOR2X1_36 ( .gnd(gnd), .vdd(vdd), .A(rst_bF_buf2), .B(_208_), .Y(_204__4_) );
	INVX1 INVX1_47 ( .gnd(gnd), .vdd(vdd), .A(d12_5_), .Y(_209_) );
	NOR2X1 NOR2X1_37 ( .gnd(gnd), .vdd(vdd), .A(rst_bF_buf1), .B(_209_), .Y(_204__5_) );
	INVX1 INVX1_48 ( .gnd(gnd), .vdd(vdd), .A(d12_6_), .Y(_210_) );
	NOR2X1 NOR2X1_38 ( .gnd(gnd), .vdd(vdd), .A(rst_bF_buf0), .B(_210_), .Y(_204__6_) );
	INVX1 INVX1_49 ( .gnd(gnd), .vdd(vdd), .A(d12_7_), .Y(_211_) );
	NOR2X1 NOR2X1_39 ( .gnd(gnd), .vdd(vdd), .A(rst_bF_buf4), .B(_211_), .Y(_204__7_) );
	DFFPOSX1 DFFPOSX1_15 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf0), .D(_204__1_), .Q(d13_1_) );
	DFFPOSX1 DFFPOSX1_16 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf4), .D(_204__2_), .Q(d13_2_) );
	DFFPOSX1 DFFPOSX1_17 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf3), .D(_204__3_), .Q(d13_3_) );
	DFFPOSX1 DFFPOSX1_18 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf2), .D(_204__4_), .Q(d13_4_) );
	DFFPOSX1 DFFPOSX1_19 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf1), .D(_204__5_), .Q(d13_5_) );
	DFFPOSX1 DFFPOSX1_20 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf0), .D(_204__6_), .Q(d13_6_) );
	DFFPOSX1 DFFPOSX1_21 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf4), .D(_204__7_), .Q(d13_7_) );
	INVX1 INVX1_50 ( .gnd(gnd), .vdd(vdd), .A(d13_1_), .Y(_213_) );
	NOR2X1 NOR2X1_40 ( .gnd(gnd), .vdd(vdd), .A(rst_bF_buf3), .B(_213_), .Y(_212__1_) );
	INVX1 INVX1_51 ( .gnd(gnd), .vdd(vdd), .A(d13_2_), .Y(_214_) );
	NOR2X1 NOR2X1_41 ( .gnd(gnd), .vdd(vdd), .A(rst_bF_buf2), .B(_214_), .Y(_212__2_) );
	INVX1 INVX1_52 ( .gnd(gnd), .vdd(vdd), .A(d13_3_), .Y(_215_) );
	NOR2X1 NOR2X1_42 ( .gnd(gnd), .vdd(vdd), .A(rst_bF_buf1), .B(_215_), .Y(_212__3_) );
	INVX1 INVX1_53 ( .gnd(gnd), .vdd(vdd), .A(d13_4_), .Y(_216_) );
	NOR2X1 NOR2X1_43 ( .gnd(gnd), .vdd(vdd), .A(rst_bF_buf0), .B(_216_), .Y(_212__4_) );
	INVX1 INVX1_54 ( .gnd(gnd), .vdd(vdd), .A(d13_5_), .Y(_217_) );
	NOR2X1 NOR2X1_44 ( .gnd(gnd), .vdd(vdd), .A(rst_bF_buf4), .B(_217_), .Y(_212__5_) );
	INVX1 INVX1_55 ( .gnd(gnd), .vdd(vdd), .A(d13_6_), .Y(_218_) );
	NOR2X1 NOR2X1_45 ( .gnd(gnd), .vdd(vdd), .A(rst_bF_buf3), .B(_218_), .Y(_212__6_) );
	INVX1 INVX1_56 ( .gnd(gnd), .vdd(vdd), .A(d13_7_), .Y(_219_) );
	NOR2X1 NOR2X1_46 ( .gnd(gnd), .vdd(vdd), .A(rst_bF_buf2), .B(_219_), .Y(_212__7_) );
	DFFPOSX1 DFFPOSX1_22 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf3), .D(_212__1_), .Q(d14_1_) );
	DFFPOSX1 DFFPOSX1_23 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf2), .D(_212__2_), .Q(d14_2_) );
	DFFPOSX1 DFFPOSX1_24 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf1), .D(_212__3_), .Q(d14_3_) );
	DFFPOSX1 DFFPOSX1_25 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf0), .D(_212__4_), .Q(d14_4_) );
	DFFPOSX1 DFFPOSX1_26 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf4), .D(_212__5_), .Q(d14_5_) );
	DFFPOSX1 DFFPOSX1_27 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf3), .D(_212__6_), .Q(d14_6_) );
	DFFPOSX1 DFFPOSX1_28 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf2), .D(_212__7_), .Q(d14_7_) );
endmodule
